`timescale 1ns/1ps

//Author: Richard Barrie

//Single part link with analog AWGN channel

module sys3 #(
    
    parameter SIGNAL_RESOLUTION = 8,
    parameter SYMBOL_SEPARATION = 48,
    
    
    //random seeds
    parameter [63:0] RANDOM_64 [3:0] = {64'h2629488426294884, 64'h588f503226294884, 64'h2629188426294884, 64'h2645841236254785},
    

    parameter M = 10)(
    
    input wire clk,
    input wire en,
    input wire rstn,
    
    
    //amount of RS FEC symbol IL
    input wire [3:0] n_interleave,
    
    //for loading markov model probabilities during reset
    input wire [63:0] probability_in,
    input wire [31:0] probability_idx,
       
	output wire [63:0] total_bits,
	output wire [63:0] total_bit_errors_pre,
	output wire [63:0] total_bit_errors_post,
	output wire [63:0] total_frames,
	output wire [63:0] total_frame_errors);
	
    //parameter [63:0] RANDOM_64 [3:0] = {64'h2629488426294884, 64'h588f503226294884, 64'h2629488426294884, 64'h2645841236454785};
    
    wire binary_data;
    wire binary_data_valid;
    
    prbs63 #(
        .SEED(RANDOM_64[0])) prbs (
        .clk(clk),
        .en(en),
        .rstn(rstn),
        .data(binary_data),
        .valid(binary_data_valid));
        
    wire [1:0] symbol;
    wire symbol_valid;
    
    grey_encode ge1(
        .clk(clk),
        .data(binary_data),
        .en(binary_data_valid),
        .rstn(rstn),
        .symbol(symbol),
        .valid(symbol_valid));
    
    
    // Generate voltage levels
    wire [SIGNAL_RESOLUTION-1:0] signal;
    wire signal_valid;
    
    pam_4_encode #(.SIGNAL_RESOLUTION(SIGNAL_RESOLUTION), .SYMBOL_SEPARATION(SYMBOL_SEPARATION)) pe(
        .clk(clk),
        .rstn(rstn),
        .symbol_in(symbol),
	    .symbol_in_valid(symbol_valid),
        .signal_out(signal),
        .signal_out_valid(signal_valid));
        
    
    wire signed [SIGNAL_RESOLUTION-1:0] noise;
    wire noise_valid;
    
//    reg [63:0] probability;
//    reg [31:0] probability_idx;
    
    random_noise #(.SIGNAL_RESOLUTION(SIGNAL_RESOLUTION),
        .RNG_SEED0(RANDOM_64[1]),
        .RNG_SEED1(RANDOM_64[2]),
        .RNG_SEED2(RANDOM_64[3])) r_noise(
        .clk(clk),
        .rstn(rstn),
        .en(en),
        .noise_out(noise),
        .valid(noise_valid),
        .probability_in(probability_in),
        .probability_idx(probability_idx)
        );
        
    wire signed [SIGNAL_RESOLUTION-1:0] ch_noise;
    wire ch_noise_valid;
        
    noise_adder #(.SIGNAL_RESOLUTION(SIGNAL_RESOLUTION)) na(
        .clk(clk),
        .rstn(rstn),
        .en(en),
        .noise_in(noise),
        .noise_in_valid(noise_valid),
        .signal_in(signal),
        .signal_in_valid(signal_valid),
        .signal_out(ch_noise),
        .valid(ch_noise_valid)
        );
        
    wire [1:0] symbol_r;
    wire symbol_r_valid;
    
    hard_slicer #(.SIGNAL_RESOLUTION(SIGNAL_RESOLUTION),
        .SYMBOL_SEPARATION(SYMBOL_SEPARATION)) slicer (
        .clk(clk),
        .rstn(rstn),
        .en(en),
        .signal_in(ch_noise),
        .signal_in_valid(ch_noise_valid),
        .symbol_out(symbol_r),
        .valid(symbol_r_valid)
        );
        
    wire binary_data_r;    
    wire binary_data_r_valid;
    
    grey_decode gd(
        .clk(clk),
        .symbol(symbol_r),
        .rstn(rstn),
        .en(symbol_r_valid),
        .data(binary_data_r),
        .valid(binary_data_r_valid));
                
    prbs63_IL_FEC_checker #(
        .SEED(RANDOM_64[0])) fec (
        .clk(clk),
        .data(binary_data_r),
        .en(binary_data_r_valid),
        .rstn(rstn),
        .n_interleave_in(n_interleave),
        .total_bits(total_bits),
        .total_bit_errors_post(total_bit_errors_post),
        .total_bit_errors_pre(total_bit_errors_pre),
        .total_frames(total_frames),
        .total_frame_errors(total_frame_errors));
		
endmodule




module parallel_sys3 #(

    //ncores should be at most 50
    parameter N_CORES =  10)
    
    (input wire clk,
    input wire en,
    input wire rstn,
    
    //input wire precode_en,
    input wire [3:0] n_interleave,
   // input wire ifec_en,
    
    //for loading markov model probabilities during reset
    input wire [63:0] probability_in,
    input wire [31:0] probability_idx,
    
	output wire [63:0] total_bits,
	output wire [63:0] total_bit_errors_pre,
	output wire [63:0] total_bit_errors_post,
	output wire [63:0] total_frames,
	output wire [63:0] total_frame_errors);
	
	//random seed values
    parameter [63:0] RANDOM_64 [512*4-1:0] = {64'h7415d4fcbce0bca4, 64'h100706f6588f5032, 64'h3338ae9426294884, 64'h3cb3d3d062ef4047, 64'h6f3964c59150e670, 64'h749b4f9cb473e2d8, 64'h41118bd6e2bf8909, 64'h1692b199b0e9861a, 64'h742735029615e72f, 64'h31b15f9f3f8b5b02, 64'hd02dbf0ef861fdc1, 64'h5b38c811b6284d30, 64'he255597ae6b4a227, 64'h24691dc9195f86a1, 64'h38c26188e2c1134f, 64'h279a6df27510da3d, 64'hf5e4bb958ff5acd4, 64'hb60cee0d5bb947c7, 64'hb4c29df4d84f66bb, 64'h1463a1bcc408dde1, 64'hfd53a014c38f4c3d, 64'h534e7a98cd6d526b, 64'h28c634b37b7e9409, 64'hea101b935677a73e, 64'h5510eab42f34f49a, 64'h14a5e7e9b2eba7b8, 64'h42ca6e744fbb2fcf, 64'h85fa41421cce9843, 64'h99c9c923333700ef, 64'h9d6eeea4b7f12755, 64'h288f6d65735f9993, 64'hb6a7f21973672ca1, 64'h1bfd23f9909d79a6, 64'haf4f8b038b92c97c, 64'hf2b3e6dd9cc5f113, 64'he8d1038130fe7222, 64'h316d2387d1c61eec, 64'h6f7143cf37af5ca4, 64'hee9a208f6376bc04, 64'hc431e548be3d50f4, 64'he3fe5385a5ae6ba0, 64'hc439e73563bc506b, 64'h50c85ea3e7033fcf, 64'h76bdec37f78fc5c3, 64'haf39d87ba534fc2d, 64'h2b89fe1af3e09ebc, 64'h7bfa99fb9ad04207, 64'h71f3ecd848e2f00b, 64'he8cfa34499aede20, 64'h10b05a58a41d622d, 64'h5e6510128e7e7327, 64'he4a0485865bea771, 64'hea0c6651a59b3edb, 64'h13cc0ea3ef109fa7, 64'hb5d0b4e5ff5b8415, 64'h395c99d130e99ed7, 64'hefd2aa4eb73c8202, 64'h1fd70cf5c54fa664, 64'hc4ee272ded86a0a2, 64'hbac414c82dd3353a, 64'h14c56f78164a672e, 64'h16cb26904b173540, 64'hde681dff9151c7d5, 64'h94ad61e4da1660c7, 64'h2dcd356053010b95, 64'h9c950cb6f8b3f679, 64'h96a5b25a1479b081, 64'hd026df1547e9f07c, 64'hd1b48b116d162871, 64'hdf4002f5c34f275b, 64'h957f666530bfcf1f, 64'h1e6157c52d1f5789, 64'h1ab1447629cc7076, 64'h462b94efbb1e0b00, 64'h965502ea1303707e, 64'h21461989f825752d, 64'h985817a740ca561b, 64'h4c8ee4cdc284a915, 64'h3ee72ff59b86b148, 64'hf8ce0734db3d295d, 64'h49903f0f86813615, 64'ha4ca1450d6f49623, 64'h35a1436714755266, 64'h20ce291884b90b2b, 64'ha184e1d398863b78, 64'h5c2abf16fd449398, 64'h9b238bd96b3bdfa8, 64'h943a4233c2e158f2, 64'hb09dab424f94a85a, 64'h1feb9cbb68d1f91f, 64'ha721d7f942711757, 64'hc4a94d1d1ff8005d, 64'h4e79c279d1241ed3, 64'h3e6c9a32a97879fe, 64'h8debbe6aedf433a3, 64'h4f30f41e1fd4a640, 64'hc06a73eac9529e3f, 64'he9e034bbefac5d2b, 64'h13592f45483f34e2, 64'ha406dcbdf3c39010, 64'hf40ad21e9598c59b, 64'hebbedaa9a9f9d3f0, 64'h6d9a12ef84a34440, 64'ha108d60993e4396c, 64'hee48963dec7efb78, 64'h6ec5285df72ed98a, 64'h39bfd60f2e51af89, 64'h306b4373895be22b, 64'h152a7beaf3834a2f, 64'hd681f97d139ac425, 64'h3a497f7a5fb1fc6c, 64'h2f707237d2471baf, 64'h62bc9eb5f1a03427, 64'h9baef383e2eb6fe8, 64'hdabc7bfde94b4dd7, 64'h7e5f0b25931f8c63, 64'hcfaa3464549290f6, 64'h85a92d2b9fc9565a, 64'h13ba5d4d9e6f7f6b, 64'h7815132cd1c43b1c, 64'h5ba8a406e64b150f, 64'h9aaf8c1d3c299638, 64'hcd1a5f44a2e3320e, 64'h1cf02f8974d8b320, 64'hb2f9fd44ec76e4ac, 64'h1018b34ffa6c1506, 64'h6a611834f9b542b7, 64'ha121c1dbd6ec4955, 64'h99ee465da6bd006b, 64'h5489ce879cd70a5b, 64'hc4015651ddfecd58, 64'hc5383feab788a32a, 64'hdf799dbf5d71853c, 64'hb0fd43697c35b1d5, 64'h6bb464a272983fd5, 64'h705ae7d65c2c11d4, 64'ha542b9d977426470, 64'hf9b66651b2ac1637, 64'h3fa8224b76688291, 64'h62673167cf6eed99, 64'he3331849e8ec0cbe, 64'haf0d815a50d9987b, 64'h4c9168ffdd2cedfb, 64'h8ea6c9b2d084c6ea, 64'h9965b1cbbff446da, 64'h8c90130cc9031b83, 64'h9886a28d7fc53707, 64'h623ece78205ec84a, 64'h6ab3a95e231c39ea, 64'hfbe048923b964b29, 64'hd2d89930e1fda4bb, 64'hb5381c3898adbc9a, 64'h36a215c8800d1bce, 64'h62d75eef4602747c, 64'h9e33ede25af1dbdd, 64'hebe9d02fea5001b5, 64'h4db559152a9d295a, 64'h3e4fa15987e67392, 64'hbedc4daf41f77760, 64'h4b872e8ddc66b852, 64'h73cdbec9a401216b, 64'h481472962878de51, 64'h8bce415082838ad1, 64'h34a42555a53bc65f, 64'h928ffb51acfe32d8, 64'h32b0e0c4c45dde7d, 64'h454ab2fc8ca4f9e1, 64'hcc789686155bfb44, 64'h5dd8d45ce18059cf, 64'hdabaf5539139ca3f, 64'hdffc6991f3f41483, 64'hd6567229dcfcda56, 64'h27b2cb6cac502360, 64'hb8d81571a275320f, 64'hcfe85c98184c0e46, 64'hc8db77c6bf9d67be, 64'h4e53de8a4db25675, 64'ha7c0b74162df1378, 64'hcf2e688c7b133979, 64'hcbdc1fc2fdb6961e, 64'h580f420c32524731, 64'he85063ed91f96883, 64'hf9f00c63a8c8f96f, 64'hfe8a0428930e9718, 64'h8e579c013080b0bc, 64'h655e8695164ade69, 64'h367eae0ac2f3f2fa, 64'h174bc1c867f8686c, 64'hdef68dc5b63e1e75, 64'hb5d37c373d45d856, 64'h7a0e99599b941dad, 64'hfd8a584d40efff9d, 64'h4b74b5a14eebea0e, 64'hc40a97d47dac906b, 64'h1da9bea58a0b3ce2, 64'h42ded520cfaa3eac, 64'h575c0a4316a01d07, 64'h9e6c7d5dda858e53, 64'h6b71a174c3f74b6c, 64'h8aac884e91d41433, 64'hf643a50bd0f35b70, 64'h17c1ede1ba40c0b2, 64'h7f99b0e8f369682f, 64'h4524d3c45018e7a7, 64'h238dc2aa76de5741, 64'h2a2a1ce5a81bdbcc, 64'hd0b60fb2b73b6c28, 64'hc7e406fb62306192, 64'hdb011d7976e78db5, 64'hd5c32a9ca65bec8b, 64'h326be98122d01755, 64'h14665b8b20039578, 64'h7e0f63b82b33ba4d, 64'h16ab024bc52ab07e, 64'h6ec39d10c343e6b4, 64'h7c93c0a87c05546a, 64'h82bcc65b81c2cd1f, 64'hd0c25b127092ff16, 64'he91feaee18e507e2, 64'hc9bad6f22e27680e, 64'ha471793b127cc7bd, 64'h914542a010b96c5b, 64'hf44958a0e94be6a5, 64'hcf08357cebaa7448, 64'h32ef190535daef7d, 64'h3d08170aa56625f3, 64'he964ef79fd96d89e, 64'hbaab5d27bfa1d130, 64'hea3af9787035aea0, 64'h4bf6d368399f8cb9, 64'h2cab70f1d306cb67, 64'h333aec664f6e6ff6, 64'hd494d6d25a8a7b13, 64'hfbc7ba644ffe4828, 64'h9013a95a5b78da6a, 64'hea95e1fc67f93d7e, 64'h780fe9a08af34355, 64'hf1552f68176d81c8, 64'hbc0d066de5d8345e, 64'h168c86eb8d4ad422, 64'h5e3cd065de47061d, 64'h960b41c4b5a799a9, 64'h7caf51ada6cb4ea9, 64'h559f8cf3123e606b, 64'h9a6be2795abf21ed, 64'h8c24ebd8ebeff9c2, 64'h765a9c6b4b600333, 64'h691c49e8efa58c09, 64'hf0d93180daa3a1ce, 64'hecd97cfe46b2319e, 64'h24fee82f468de903, 64'h5b734c9f39f19d8e, 64'ha1b3dd867342bfd5, 64'hd3eca30c3c6e6964, 64'hb8734b4349af7319, 64'h99d0055563c1cc48, 64'h1dabe48946ea4fdc, 64'haf62760587570bb6, 64'h8c90579239eece58, 64'h98f8c82cff3887cc, 64'hd40a595e9ea64107, 64'hfa3cc4b4e8600155, 64'h9ef226c517c84600, 64'h267560741fb0702d, 64'h7c6a7c136a1ab756, 64'hfa1581913850e4bf, 64'hf97811d5c831a7ec, 64'hd5d12c41a7d3ea71, 64'hb07ef1008273a68c, 64'h1327190864b8b1a4, 64'h8618e439bf38cdd4, 64'h807886807dc6f543, 64'h3109ffb2129d00fa, 64'hc5fc9dc85cc9e702, 64'hfc4084e944db30dc, 64'h614a389a8dbc2db8, 64'hc52c87f87f536c19, 64'h2df518d95b0015af, 64'h8915a865b1b94877, 64'hc8d603692f47d494, 64'h157fe7da8c946afa, 64'hd265b4d61306601e, 64'hb1648c19b4d57f59, 64'h7bd1b876eb8c9def, 64'haaa58b891141ef86, 64'h844348a1de3c7c6b, 64'hd74bbfe5abcc08ac, 64'hb1b007fb9ad703a2, 64'h51c9eb439686f66f, 64'hb13713f7649546c8, 64'hdd66184b3ecf1a68, 64'hc35b63fe55813157, 64'hc9b63a6c76a82e78, 64'hd1d8fd8264d92e96, 64'h43495002c825f5d0, 64'h5a12f616bffa93b4, 64'hc2ac6e3745229d02, 64'h43630cb93fbf5c45, 64'h323453a16a7ff475, 64'h1664046a2a9ef28e, 64'hb1e536b0cff2453b, 64'h2353bbf2479bca3b, 64'h41d4854bec28f960, 64'hbab729fc94eeaba7, 64'h591595cfd85d6ec5, 64'h787932b3eda1265e, 64'hb973d2a782ba3e5b, 64'h2e4a594afa401da2, 64'h365c2df3409fdfe5, 64'h777bce9a71022a44, 64'h33386936bf095abb, 64'h3d4c7f36aa88f2ca, 64'hc5088ec0429365ef, 64'ha03aa107c3be28cd, 64'ha92c28589f4f8062, 64'h56ea6e80bf95e6cf, 64'hf2dfc02576227de8, 64'hcbb940371d794e34, 64'hd87716573e23d74e, 64'h6ed2c06b5804fabe, 64'h23399161e91c8761, 64'h68d645ce8f5e0cf6, 64'h869680de2fb7fb07, 64'h418c899222490a5a, 64'h89e6b5924ec59abf, 64'h65b1dd8229ef88a7, 64'hcd032f5f2994836e, 64'hfc91f33c3a84c82e, 64'h996091f31ac34c20, 64'hcce86cc33d8163b2, 64'h8eb26ba2c19e5d40, 64'h33fbca5a9442cbc6, 64'h43fcf617c635015a, 64'hbd7fe8d53a5f2c34, 64'hdedf39ae14befb6c, 64'hde74f60d96230cd8, 64'h70c5dda6c6196955, 64'hbc101e2dfcf551f8, 64'h52bd8b9f10e9154f, 64'hf022f9ecdde532b7, 64'hbeec99118c015bdc, 64'hb9ab6447cb53bc69, 64'h69f860c3c8e09db0, 64'hc4265bb2a32bb264, 64'h7072a473b75a9ace, 64'h10bf4106c9f9a665, 64'he723d608496f8e9c, 64'h2cfbef9144de3f8b, 64'h5880d2bce3ed4586, 64'h925c253e54cf9053, 64'h3134831c55a279cf, 64'ha3543d615dcb1240, 64'h7dc435a67a968e19, 64'hd6c0a2f67652d4a2, 64'h62f7bc4fb1fe4162, 64'h4527db868023955c, 64'h5b8b342fa672021a, 64'he291070f7b72031e, 64'hcc4510567dabf900, 64'had7ebaeb2fa44f3c, 64'h77ea6240ea3c20eb, 64'ha150a13dc806a172, 64'h8920ce2d878889a0, 64'hda4bc42520460edd, 64'h9995d92ff2435528, 64'h8c4952453eabfab6, 64'hdb8165734c64b57b, 64'hb82c9b9291a9a1d7, 64'hf3b88066a5d73f3c, 64'hd91d5db211e7655b, 64'hfd710d9522a6c880, 64'h5d4fa328f3139a6a, 64'h122537edd5748813, 64'hdeb0d7d3798f348a, 64'h4d60fc16d0a53e7d, 64'h82afd770303dc39e, 64'heeaf0ac9e7086510, 64'h85f888b6dd9bcd28, 64'h74756f15b408155f, 64'h6f848b7e8960ca21, 64'h3d7e0e7ff798eb65, 64'h569c9ca528d48e1d, 64'h32a2bcfb1361d4a0, 64'hbbd3b42b977ac6dd, 64'hceb2e4d789b2fd91, 64'hce097c14b6fbc0da, 64'hcaaf02ab718e4eb7, 64'hab7707183b268fc9, 64'h5d3c9e5a396cd3ef, 64'h7212abce49f0c494, 64'h71a9498efa0da925, 64'h5ce06b5dfbcc3e61, 64'ha8b6a5fc6a059799, 64'hddcbd8fea4b368c6, 64'h4c7ce996ce490d88, 64'h77e7bdf365cd7c73, 64'h5f443709b75e57fe, 64'h5079dd16d1fc99e6, 64'h56de8b259296d15c, 64'h8519e57fdd491916, 64'he53676693c409484, 64'h9c7bcf30e791b7d1, 64'h7b117123ed3f96b5, 64'h52f53348a21e965d, 64'hb3c9f4b846c4f5d4, 64'h134de0407403852f, 64'hf13c53d36253a5a7, 64'hcb237d5139efcc90, 64'h6211951032b4157f, 64'hbc06661ab7d575dd, 64'hb53d46754cd0a701, 64'hb62a9b1b468d2932, 64'h75ea71136942e529, 64'h65461e3c1dd64fb6, 64'ha7985e67b9c18836, 64'ha342e3b0ab9855f3, 64'h38c9285133de02e7, 64'h8b66ea29e2147156, 64'h3c2619767f14d5e1, 64'h76f19a4587597295, 64'h36c338c4622f8d91, 64'h4ed9ee9adaafbc43, 64'hd01469c77664b5bb, 64'ha1af07a932e96838, 64'h8a4ea40c57446dd0, 64'hde50f460b12f0129, 64'ha808a4b22df0b84a, 64'h80f0eb59fcc70816, 64'hf3978053aad20fcf, 64'h3469f9e1a963f41f, 64'h97c247bb807ad43e, 64'h76ba9f449fd32240, 64'hdbfe2664c444e071, 64'h9b0be95fededd32e, 64'h1f899fe5fdec545a, 64'h1cb7fc163fe101a1, 64'h7575ec6d29cd586a, 64'ha5ae4f601b84a9c4, 64'h544f4a901ea617fc, 64'hb8d83a4bb06df26b, 64'h6adbfddd3d2aa7c5, 64'hc347fa0961b0e754, 64'hcedf4dc18518a23b, 64'h8e29217316d67a51, 64'haa9d9d85642855e4, 64'h47025b5d7821cb6e, 64'h6bcaccf380bfd6b0, 64'hfb1375116773637f, 64'hc9dbc23494aa0a88, 64'he56436d165304d9d, 64'h4aecaaf0eaa505a8, 64'h1a72bec4f42e4a67, 64'h9589a4126a53c18c, 64'hfed003c31e01cd0d, 64'h8c02705217769ab5, 64'h991509953b4ffc36, 64'ha76e221efb6bf35e, 64'he1fa03447c70d1b5, 64'hba07d5fbca97ae15, 64'h86c328bb8ed918ff, 64'h3430318668a7ee73, 64'h322212e4be745a2b, 64'h827badab7bbb1da1, 64'he4a3b7228ea0e5bb, 64'h722e8a6d5088b9d1, 64'h21486b61745a48b8, 64'h162e4b4155e07f84, 64'h88d79fd2f7d2ed72, 64'h2a407c7bb187a473, 64'h87fbd84bca80ea4b, 64'h327736c623f7f851, 64'h6fcffdbacf455c5b, 64'h3e008eb2c8443b0f, 64'h55abe8b1440dd021, 64'h1403017c6fad9cd7, 64'h6b75a597ae3e2724, 64'h210539fe349ffd2d, 64'h13fa6c192b4fa5ed, 64'hac6deee170a33cac, 64'h5d0bdb5495e61ce9, 64'hfe6e35fbd846d9f7, 64'hb7e8d92cec61cec7, 64'h1988ee8720e14963, 64'h81c2f24b63ccd88a, 64'hf0f0c447857edf08, 64'h91840a95e6dccc00, 64'h7b3141d9e27cfe2e, 64'h4cdc100c51b6de44, 64'h5ece8619936a594a, 64'h44d4b4abb1249bb8, 64'h3245382426958558, 64'he0d894b648d93691, 64'h6ca41621992b8bd3, 64'h8e3145e6223ee83c, 64'he1ca4c28f445c5bc, 64'hd30072e3541cc8e5, 64'h8eaee83c6175c377, 64'h951ec274f9db5961, 64'h5acf06fbb082dd0d, 64'h5e3b6cdcc9dfe21b, 64'h5e31c3ade58efdeb, 64'hc468ec21c7081daf, 64'h80accaa142955efc, 64'h19f43a995d3d2957, 64'h18e833beb68679fb, 64'hb0e24e5477502fb4, 64'hc844f46d90a45ca7, 64'h1990fe703059b06e, 64'h3e6b80ea608f2f17, 64'h1c8e1b81a13a6000, 64'h8ae50790a430cdf9, 64'h77c3ed81db72b77f, 64'h7cf9636f13b2646b, 64'he1894e9bad7d05ea, 64'hd5854e8cf46d193d, 64'h1c380e8e486ad0ba, 64'h1f33d2387532a918, 64'hdf51a9a72396fa3e, 64'h818bff972e215e61, 64'hc97e1766d9f0fa32, 64'h1a63cb9584beeb55, 64'h49756a21f497fd39, 64'hf288c358a3581ae9, 64'hf9a310d262c447ed, 64'he77bf2b7784d83e2, 64'h48987389f1cc7856, 64'hb4365b681f942af6, 64'he0e6e739b854ce29, 64'ha12eb503bfc51d23, 64'h4cd34b77a01e0a9a, 64'hd38233d71cfcbe49, 64'h2f52935eda2fdede, 64'ha4672b938f8252b6, 64'h4b96fb7e56d1a0af, 64'he171d686753327b1, 64'h1f76984ce746c33f, 64'h40cfb7e8d64b6b77, 64'he39ffcb284d1f73d, 64'h9fa1abb68e8b5002, 64'ha5f50534dd35c36c, 64'h53b6a5d1e419f03d, 64'h983ee4d62b9fee4c, 64'h467af39c9f092864, 64'h497793a92f8a2d9e, 64'h36d7ec6fdac4f7b0, 64'ha08629e8f7418fd5, 64'h62f687e79ef334bf, 64'h9fc1a7faa3c4df15, 64'h1e33d8fdc4137ce2, 64'hf391fdd89052ae68, 64'h3e36a456c4b3c4aa, 64'h11c1ad705ec80e16, 64'hec39bbe89d3549f8, 64'hdd3ee41ca11f0d08, 64'hd56b33a3e31377ba, 64'h5d0967222d825757, 64'hbd1ce0a279aeecce, 64'h2e6aa4599d8ec3d4, 64'h18a8098a400b3072, 64'hcd3139a012e73996, 64'h58cd8ede152156cc, 64'hff657a5c9bafebf8, 64'h566909dfeef2a7ab, 64'h89b56ada7d204a5c, 64'h9d16d34a4f649deb, 64'h5944e9c26932750b, 64'h4aaae2959c4a9584, 64'hb700c95721446fed, 64'hf90f5bf2c4bca93e, 64'hd17aaa2cc464c954, 64'h2336f24b839b6b6d, 64'h7af6257eb164b83b, 64'h7bb26acdb90903e4, 64'hb3984a20b750ce3d, 64'ha476d463343c419a, 64'hc697b3f3cb737490, 64'he8fc1664481abf9c, 64'h3a6726b56ddd2150, 64'h5cef7e0bd3b6e70c, 64'ha33f0802c66681f7, 64'h76a3be6527dda0d1, 64'h2b9bc04b699e225a, 64'h3e8601c0d4faaa36, 64'h9fe9a2e9b552a719, 64'h85ddcbc925296417, 64'h486b2b857ec8d4f5, 64'h3fa97643161d428b, 64'hbf0e31d1bdfae28d, 64'h5f4b44d7da704774, 64'h76d38178df865116, 64'hadb219869b72d4af, 64'h402cb2668f175800, 64'he6a9ed845932d473, 64'he106e5f3ea194f40, 64'h5f29a662b3f016ce, 64'he7d02299222ad101, 64'he2dc70363dcd2ba5, 64'hdbf1cd45b01bc744, 64'h62a4333f345483d9, 64'ha87d311fdb7818f0, 64'hd53e6cf4a6c70a75, 64'hf5832a2e9d94e07f, 64'h3f7ad8a7770a1461, 64'h60d1ac96fe1119fe, 64'h6b41baf7fe3f8aac, 64'h8c83554b3958dd68, 64'h21e5d4b968df94f3, 64'h2d9edad1a848d477, 64'h73573c3ffdd1db42, 64'hef30793933d10fd4, 64'h6ec590f47ec7751b, 64'h96a0b108cb4988ee, 64'h84ed319c74cc6762, 64'h4ee1430aea97ede0, 64'h15585c97d511babc, 64'h3d3b7f9db494e766, 64'h6540109df9cf9fb6, 64'h2d771ea13d044b51, 64'he57758809c047be6, 64'h5a38190f102ef6bf, 64'h469f9ae532e5996b, 64'h40d2f964e71e0ed2, 64'he18aeb2ab811c876, 64'h80eb6092d6833c6a, 64'h86ff92e7673cbea5, 64'h52250dfdedf0135a, 64'h6ce09e5a864a99d3, 64'h4d10ad51e46457ca, 64'h6bfbb4f0576afd92, 64'hbc3908d43dcf0ca0, 64'h2c5dc152d8e124cd, 64'hc297b6059db9951c, 64'h4a4b4225a5944dfb, 64'ha9348d095e9ddddd, 64'h20328b95e3544a9c, 64'h7e63bdd7c75456fe, 64'h4ceeeab99deed418, 64'h76e92cb66bb44374, 64'h2e6945334a9fbe69, 64'h230abf3358af9d3f, 64'hc20257cba39a90ef, 64'hb160f01c12030e71, 64'hb2cf7b2f88c36bf0, 64'h476b03e439f9a43b, 64'h3c655a79da9f55b0, 64'hfbd25111eb4c299d, 64'h635e6090cb40ff89, 64'h93262b89d3f2388e, 64'h84182f139d969b97, 64'hccf1775a280e6a9e, 64'h90e1b79f67d6044f, 64'ha1089cccf61cd39a, 64'h6e470ab06e5042d1, 64'hcdc0bca5aad19dea, 64'h6e883bc3b55965ef, 64'h70f5dbdf30aacace, 64'h7c2785be6042ba3d, 64'h445002d6ee2f9a94, 64'hb58371d79fb78e37, 64'hc332a2969212b3b9, 64'hb820c082ef559866, 64'hdf072b73382fa0b3, 64'h4f2742fb212fbc4f, 64'hfae1a83b48bb7064, 64'hae8b29ba2582e900, 64'h4295c44688ad87b7, 64'h29305a786d5461c2, 64'h911df72d6168b483, 64'h956a824c90d30bb4, 64'h6dbf1bebb71ad57b, 64'hb2d5f644b4f3e7cf, 64'h96c205e065f06e10, 64'ha3259f34f093a2e0, 64'h9f40d4bbfb1a0534, 64'h79d7725fc181c24d, 64'h190661dfc788ce01, 64'h8c6338661146a5d6, 64'h52872ca8905c17a6, 64'hc84fa3a61cbe0253, 64'h93c5d7f6d03d1b03, 64'habe66206ef8c1ac8, 64'h21ef7fff526efd34, 64'hec9df3c8c799ea94, 64'h9ff00bf9d7e99011, 64'he70ce981f973f041, 64'hffa5199731840e19, 64'h20ee1a6e21a1ca8f, 64'h1389dbc8f93ca013, 64'h26be7ab7da044f84, 64'hb47107688503832b, 64'h6334eefb64e01ebb, 64'h4cebdc67eaa4f1be, 64'hbe277a5e1638e177, 64'h7ec3dda653832673, 64'h16f3aeb7e452db08, 64'hc90a91b75f22ec5c, 64'hcf2c8f445de9c74d, 64'h59e44c20eebf0594, 64'hfa75baa08da73ce9, 64'hf476e58ee51e812d, 64'h8c53ebac6975afb8, 64'hba7c2f707d5abb66, 64'ha14047c1fdb28e87, 64'hc9bd6a166039f13d, 64'h255c0cfa3c609977, 64'h8e71c77e741ac5c8, 64'hd0288787eff7f3a0, 64'h3ab00297de6a809e, 64'hf5c65823f645dfc5, 64'h191647041dd1ee3b, 64'h1164311c5b0b2158, 64'h1d5e1c495686e93f, 64'h6571a725f4e1ea80, 64'h8277dd5c52c6f84c, 64'h88b8a3a2aa67e931, 64'h2ab2ef23c5ef4eec, 64'hdc778c57da9eb61d, 64'he5b8bd636ba46599, 64'h7a83643228612a78, 64'h463193cbf91dedfd, 64'h544f4bf2e9c66b43, 64'he5bb8851ed66ad23, 64'h3579d44ae32220e6, 64'ha7adc50f428cfecb, 64'h62d3ebfc3661690f, 64'h7aa4c035241b2218, 64'h37ad2b063f53be58, 64'hb5d8b84a99b672c3, 64'he198f92e4ab65127, 64'ha71b1ce5184374fb, 64'h8be33bc4df2ca292, 64'hfc30bc20125e987a, 64'h4cae94a745b952e1, 64'h1b68b5b51270fee8, 64'h85a599991aea6c4c, 64'h52cc7af9a998099c, 64'h56b9e10950b795b9, 64'h9dbb2da76b540383, 64'hb89b03e58711db07, 64'ha7f8609764d08c77, 64'h54e3fae52ff83ebd, 64'hf0e63807d1291d48, 64'hf12079443c7dc78a, 64'heff5170ff094ad56, 64'h540cf99551e9873a, 64'h9457f4b53c782bbe, 64'h7a1ab1373c79ea8a, 64'hf35ec6c386849643, 64'hf7571b8eaac93764, 64'h843c5c71f83f3228, 64'h325d9488a7c258f6, 64'haeda6bdc781f1e76, 64'h1e3ee86e8640e06a, 64'h7fa1d45ad19e8629, 64'h4d9940516df17b44, 64'h49a42e30b4bf155c, 64'hfd92707b3a954550, 64'hd525b00f476fefe5, 64'h1dea08b33150e30a, 64'hf06fceb4e54006df, 64'h556c2a34f3769fcd, 64'hdbfbbb6a785130c8, 64'h8054f6f4a72a2b6e, 64'h35ed79d8138c361f, 64'h4fb90ef113b4db54, 64'hb1e13581945a3ecb, 64'h5d320fe4cb3fa1b1, 64'h32fd0e914ac57769, 64'h5627c1ef3f060f0e, 64'h251af3e7e0cb5626, 64'h252a4f76b41729bd, 64'h2ce56e0d129158c5, 64'h95be8f60e9b4c7c6, 64'hde827528613a73fb, 64'h1684a374d034cc7d, 64'hd16fb6d9e06fe8ed, 64'hb0b7164cd1ddeeed, 64'he7664b637ceb4fea, 64'h95e0c9638978b252, 64'hb6137db9b3e5cc47, 64'h8ce011ded6d51541, 64'h896315e5d5f74f61, 64'h53a48fee3ad6b8f9, 64'hf8c4d90dc210c3b3, 64'h4e599a059b7f1975, 64'hf543501823618526, 64'h240c5779a497a4e0, 64'h45e0e11dc7a4e6fe, 64'h985b4ad1afe298a5, 64'h29e01609243a59c7, 64'ha607703e7255e381, 64'h24f0cb8a690e2b36, 64'hb1508d733d803ff8, 64'he6f998b0f3f68fe8, 64'hf6c7045bbf3845b9, 64'h71825c6bc27ff35d, 64'h551de9f35b75cb4e, 64'ha16a45bf9ec3686b, 64'he2e0ee2e4d1aaba2, 64'hc7e29cf8f1d7dae9, 64'h103f76a18242ea59, 64'hadb08ecdda65c73d, 64'h3c18f311dd7a6c70, 64'h67729d77e6254f6b, 64'h16a69bfc247e5ec3, 64'hfb89dbe9a247cc5f, 64'h743b54d6389c84ff, 64'habf9ed4618dfbf8b, 64'h5ac98f115da28fd7, 64'ha1c93adeac33128a, 64'hdb0d9837ee9e92b8, 64'hae8285d69ac3016c, 64'h6fb11540f7fcabeb, 64'h34fa9fd4e6d2222f, 64'h5aa4a49593a32b70, 64'hb3b226a348c0b205, 64'h3841bdf08a09228a, 64'hce0c1dd4b62df1cf, 64'h2c8db8cbe82d9a09, 64'h8323137df333d0b0, 64'h94d2f788245a3954, 64'h40975434dd04618d, 64'hb96c2d6ce6c91589, 64'h5efebaf98eb867e4, 64'hac1876169ea13ae5, 64'h478d1530766fe75a, 64'h4b8bf7e6daf29552, 64'hfccd76541ffa1c33, 64'hbb57bd025f3a4cae, 64'ha61abfe94df37c54, 64'hac3de85369134874, 64'h56c1cb7bead2baba, 64'hf233217fa340837e, 64'h4378e685f175e53b, 64'hc41bddadc442f530, 64'h42d028a8d73cd125, 64'h499f723fa796c752, 64'hba93d6d5c22c09b6, 64'h6da9dd0cc65bac21, 64'he8b461c09cfb1603, 64'h25b2c5df2ef448d3, 64'h2943546439746017, 64'h2e57e9f6cacace83, 64'h1975717d49f95963, 64'he2f9d6f7f9a4ffb2, 64'ha14d20cffa4c1438, 64'h1a6da9a9f3a84f97, 64'h5ab60804cfc0e42e, 64'hd28d0d58de665040, 64'h7e0d5ca1ef5aca9d, 64'h4de4f1eaf04454c1, 64'ha496b5d5fc81bc4f, 64'h17d5a39ebe0a3d52, 64'h97bba6f9862e8892, 64'h4e365c955e707a2f, 64'h4bdef53f449fd207, 64'hcfeb297088932630, 64'h23f72fd0ca79e8a5, 64'h90136635c173fc54, 64'h8bb1c9dc6ffcad76, 64'hfcb3009816c73a02, 64'hefdd03b7ef67baaf, 64'h6dd20baf4378b8c1, 64'ha49c770c3ab69ecc, 64'hd0c51c894cf1b234, 64'h55cb2153ebd1ddbc, 64'he8b335d3907dcd50, 64'hdf14d3b5649b99dd, 64'hff7e02937815e5c9, 64'h56c1400119fa5229, 64'hfd8798627f92b230, 64'hc04ce73da9cb386e, 64'hbd8adbc61c444102, 64'heccf96f8ee711fdb, 64'h947a9311f756fe01, 64'h536de880a083e387, 64'h6f26aaeda6b9bf53, 64'h5826d90ad4a56111, 64'h20bfa6891a0cf53b, 64'h1bdae9f4341bf4fb, 64'h6ee25547f54b2934, 64'h2a974596ab69a7cc, 64'h8ea110c464c736a3, 64'h3f915c5444f14ce7, 64'h1a8464c1bb28cb66, 64'hacebf11d7a813751, 64'hbc8ba4642a64ec7b, 64'hf14ae7f1db6e2f5e, 64'hae2b26a46aeb6313, 64'h73f9dc1e83b78978, 64'hf077d5b8df4326b2, 64'h82b3a42c95159dd6, 64'he218d035f3d2ce8c, 64'ha96782ecc3a516a6, 64'h6463d592ec53a8f1, 64'hd8d20bc3947e5038, 64'he03b0409dbf820df, 64'hd204cb342f5dc463, 64'h90a3ff8ae8301d55, 64'hc8ffe85e74f89e74, 64'hfab0f8ac4c2f80b4, 64'h60110331f5021445, 64'hd2177893e814e3cf, 64'h12c8107b6b24ba0e, 64'h4886781257063fe5, 64'hc11e717dbdc7c5db, 64'h7ed4f4ad67aa7681, 64'h9c5373e590170124, 64'h94239bada3b6e948, 64'h6ef4a13ec9366231, 64'h4c49ec71ad61f10c, 64'hf67ecd0110da678d, 64'hbd9b4d762a28a7a7, 64'h92824db2a675b857, 64'h4a4eabe2eb529155, 64'ha55ae1bc479b5265, 64'hc8d4ebef29525ae1, 64'h95410b2826ca19d7, 64'h9b6fa9544cb7191f, 64'habdf3d9ebbcc6872, 64'h8dcdf6d4adce1d84, 64'hd330c61cd1cd8dd1, 64'ha4b942f87c43bc3b, 64'h71e87285e1f07e68, 64'hb8b420293c626864, 64'h97c69546ea1d2a5f, 64'h342a64a4daec9b22, 64'hd4d93d5287d7846c, 64'h190526df33668dcf, 64'hed6eebe11a98dee5, 64'h69665300a491cb90, 64'h3f447ccefb758a51, 64'h356f1e4b9185e3c7, 64'ha4529da3477005c0, 64'h7fea063985d79065, 64'hc80c0640a83a359f, 64'h80364678b010f32a, 64'h7ccf82548e2bb85e, 64'hae0e6ba53b7ca4ef, 64'hcd21c3b2a0b00bdd, 64'hfb47a708455f3932, 64'h7fe76985e6f43b7c, 64'ha0581196be3ae958, 64'h7347e518b43bfbb1, 64'hf30d9efd400b6e90, 64'hd1c48596f8b06a5c, 64'h137f1a5743a67a1d, 64'h2c2ba353c82e803d, 64'h237df272ff9e8770, 64'h6d81c324e93fa86f, 64'h3d42353d79cf301e, 64'hdac13cf99edd6016, 64'h7eeafe548b093351, 64'h99bb86db79ad364e, 64'h3e74432b2b5a0e70, 64'h344b71a11c990b7a, 64'h96151426db73faa7, 64'h66304acd2213199b, 64'h762c8204a07b5c92, 64'h7618c9f7d292b66d, 64'hf20d7db0e0c75163, 64'hb8f5baac80df2a7b, 64'hb3d8f7bf13386bc7, 64'hfbcb74a3394c6e68, 64'he980a384d1b4d516, 64'hd008950c508b6e70, 64'h4498cf5176e983bc, 64'hdbd95c467c175343, 64'hf080363964a49e2d, 64'ha4a77465fb5e2618, 64'haa6e565e1aeb6910, 64'h7f40f29b60571f60, 64'h8fb93bfe5456ce9c, 64'h2d57bae1b063acec, 64'hb386be4ce01d09e2, 64'h2fc584dbcfab3b54, 64'hd66cabdaab2c072f, 64'h412e6aa94ebdb04f, 64'h747071c992082292, 64'h8295c9ba8030bc5c, 64'hd98fd031e0d316de, 64'hd4055d14e2ac1e82, 64'h990ac741f75e614a, 64'ha19215b3a0f28c9a, 64'h5ca1a729b37d2f61, 64'h1c78c59c304a8839, 64'h2f42142bad3f912d, 64'h3a146f3861e00f92, 64'h1aa282164818a39c, 64'hf769f1498a318660, 64'h344204b78d85a4ea, 64'hf2713770dfc3bfab, 64'h6e1886e95420d1f8, 64'hc6d0aeca49b75b5f, 64'h4d04092f242e43ff, 64'hdf6503607b7ee8cd, 64'h96d425dac0cf8571, 64'hcf2846a87b66e66b, 64'h3c30cc0cd6e558ae, 64'h177083c1f336fc22, 64'h9a7984d6e217e254, 64'ha20e42ad4c65f701, 64'h571238f68fe6c315, 64'hf6e615dd3c4768f2, 64'h8a60280762825751, 64'hc8bbecdad0b01def, 64'h75e4f5fd40fd4952, 64'h2019f9f93facf30a, 64'h51604ee99fb59754, 64'he18a40052ec68247, 64'hf5f71dc6b3f60443, 64'hc212485cfbe4320c, 64'h73dd3b428f947cf8, 64'hb302d7fb8b170c7c, 64'h57c97664294ad595, 64'h54623b25c88651aa, 64'ha9c9b07ad051c227, 64'h8c1be2b047b439b1, 64'ha6b5fb1658f618ea, 64'h17163f00e8ccaae2, 64'h74e3819e764579a4, 64'hc1e681b2f3a148cc, 64'h21675aa33972c13f, 64'h5d5da4e64b9f2f8a, 64'h86eb3630d5decc6a, 64'hdcf410b09effcaa9, 64'h49a446333cc21c5c, 64'hc269e9c048ee6e84, 64'h917a5202c3d3cfc3, 64'h46c7a00039e15a5c, 64'h19895c50336aa120, 64'hdc58680d291cd497, 64'h45acc06917dc9a34, 64'hb2535a08479bd74d, 64'h7343133d316ea9fa, 64'h6a883aec75dd701c, 64'h8182f776757b66a8, 64'h28a95d01c96b54e3, 64'h30edefd675d48603, 64'h5144fbca583ded93, 64'hb16188438c44d0fa, 64'h3d9ef2ca80979eb8, 64'h617d6418b9144ed0, 64'h46434a0cdacc1238, 64'h8e4b8cf58826110b, 64'h4ce274bb3cad6784, 64'h813c902ffba34ad0, 64'h2fe5c25e5407ee8e, 64'hd02764cdaf8be485, 64'h52e6eaa95b83f2f0, 64'h74c99eeaa0ab37fb, 64'hbca42c82ddc08852, 64'hb3777d1f48e02d95, 64'hee2c450bcb7ca53b, 64'h59c584a6593116cb, 64'he37afb432e424308, 64'ha807d56b52a6ab98, 64'hd6873020677c5215, 64'hc002034a3e2e27bb, 64'h838c0934d0dcda96, 64'h6f46f4ab36c71be8, 64'habc177c0c4cc5668, 64'h533f09187c53ac3a, 64'he81b94c9e146cc15, 64'hb9b99b549dd0eecf, 64'hd42bf77ae9d5afe3, 64'h109a10816f55ac89, 64'h96bd02cfc0243ccd, 64'h24fe53976ff0f24b, 64'h531becdf75a4752a, 64'h8783cea5ae6755d9, 64'h8718bf96a4e990f6, 64'h9bc91ae976ccbe17, 64'h1131bf733eaf16a6, 64'h5cd97f3133465608, 64'h9fade8ada2c28721, 64'h8805bad95d00f4df, 64'hacc82cbb3dab0466, 64'h116953d8c062d66f, 64'h7a70e045b77b6430, 64'h3c69103c1f075c53, 64'h6abefdd8b70a068e, 64'h28ad29173f000e2a, 64'h7cf2d9d1a51367fe, 64'hc407a2412a561ea6, 64'ha5e8dfdb6cf76e34, 64'hb0d25a2e40dabfe7, 64'h8eb354b83951aada, 64'h147bc2d284de3920, 64'h3c33e1f2a933d070, 64'h90c7282bc9fca4e7, 64'h6e4f74d8fd77f05d, 64'h8ba6ca7b82eae8e7, 64'hc3ddbed39971f800, 64'h66fdde7e856b331b, 64'h3d64a9696e75c3d6, 64'h1730d99f7f01c915, 64'h51dfb0838e696c27, 64'h17067aa9953887ec, 64'h5651ca3c9a990707, 64'hbfdd613a79ae5b28, 64'haf285aef4956a0ad, 64'hffa9ed924a4a74d5, 64'hf1cc7f6f4421fb42, 64'h876a5b16d5151cdc, 64'hbbfb2b6bb956dc4c, 64'h79b4ab03c5008379, 64'hecc9f2a279eca6b8, 64'h8eb633091fd939ee, 64'h6dc9190080232335, 64'he6d542ce2a88a62e, 64'hbf79182792e9bfa4, 64'ha19189701725dd35, 64'h333828b65427edec, 64'h112b56b1b0990e1b, 64'he0dca5fd9345bba1, 64'h925bffc4a3c63379, 64'h5886080968040351, 64'h99fc4bfed2364454, 64'h406218e45e9b13f8, 64'hc24d14e661d223df, 64'h1b6d3729358691d8, 64'h3e870e9786d3b41d, 64'ha86e13dfe340b725, 64'he89bd89659b7f527, 64'hc4cfabf553c860d2, 64'h68755ce656411eb7, 64'h734928aa438821e2, 64'h5c8e80102d42c0dd, 64'hf71fd73588f4b753, 64'hed8b4e52c314143d, 64'h7dd969b3c51bfd52, 64'ha6b9bceb58e6eb0f, 64'h8d32bf8cbaf47618, 64'h594676a013016732, 64'h50621178cf380ac2, 64'hef32c680a614589e, 64'h2fdfb11ec5d11f75, 64'h8e751081c4edb73d, 64'hde111a61f368f3f2, 64'had16c940dd059fda, 64'hc2389c3bbe8118d7, 64'hde1c1aa5ed854e8d, 64'he87f8caf6efae565, 64'h242a4477d719025f, 64'h9157f463921928b1, 64'hd60ac5b717ad1bb9, 64'he2b5e35d184fe9be, 64'hb65ddfa99cff0be2, 64'haa0511d669c77c9b, 64'h521c630e8a421031, 64'he498f8ea97ab65b9, 64'haf27de2f79ee5707, 64'hf95039bcc2349459, 64'h652d35d5acd8f258, 64'h923a5a34e42c69e8, 64'h5203522729efaa92, 64'h3de7c13f6ce41edc, 64'hdcf96f0e5100b626, 64'ha6537c21a5a705cd, 64'h71ee6a7f1c149723, 64'hc2c297da56f96079, 64'h6fa145886a89995a, 64'haf43bee624b85131, 64'h93f93c9a13b3844b, 64'hfbedea489f9f5e59, 64'h6c2ffa6a33383160, 64'hb7403453e964de7f, 64'h5c589a0cc7f54702, 64'h54ffe226f5bbecd0, 64'hb88e47ada600f543, 64'hef60578e5091f6db, 64'hedaaf393b2bd6a5d, 64'hc92083309931466c, 64'hd8231a78b7966f0b, 64'h332fa37ea2fd9c9c, 64'h53097101ebcf96b9, 64'h3f93645554926be6, 64'h1b6fe7b37b6b433b, 64'h95d2320499a797ca, 64'he94a62e063611caf, 64'h7b6824c6dc4c0ac0, 64'h9a706474acf55370, 64'h52ce65b384fe3c9e, 64'ha50750903003baae, 64'h17e5e95c2b37f8d0, 64'h8297356315c433dd, 64'ha64a46d0276b79df, 64'h4c3b13af765bba03, 64'h2bcc653450eeb6ea, 64'h150f2296fc6932e6, 64'ha2c7151e6ace0f53, 64'h165de6e36d8fb155, 64'h7c9d33b7ef70d613, 64'h52d74bdca38c330c, 64'hafa3f1973ca17126, 64'h896219a5ccc29b5c, 64'h272dd0dea172cf09, 64'h16411f4d11b0f362, 64'h1e49700983893e85, 64'hee2b42ad71557219, 64'h22020160deb97efc, 64'h8ca1a4c75c8b6b78, 64'hf720b4f8f12ecd96, 64'h4e6790ce405583f8, 64'h9d568cfdda34519e, 64'h60d024ce9cbe3942, 64'h36f055313eb3d6cf, 64'hc6b86f8934060caa, 64'h4fd15420b57a907d, 64'h139f164a17ba0631, 64'h5501980160ca20d3, 64'h66ee8ebad1b9c9fa, 64'h18a2abb06603cdc8, 64'ha92fcefb32522c29, 64'hdddb75e2aaef7a2d, 64'h2baba0c941f18140, 64'hc2eb6ade70d14da2, 64'h8445d72ee4fd3d71, 64'h30fc881df773108f, 64'h1a3b2aec27dd9c03, 64'h4593c4ebd1949664, 64'h7d68d346acc7c00c, 64'h39d64a6b38036544, 64'h8d00ec0cc1aba416, 64'h7efe6e60e0b516e3, 64'hae7fb5934bc81855, 64'h4860647869c56e28, 64'hc5967d92f11ae3de, 64'hdedb812e4ec95dfb, 64'h72f26ad7a2c544fd, 64'h933d824c6d6d0d7b, 64'h28574ae4baf0521f, 64'h25270644dfdbcc1a, 64'hdf3a45aeba073776, 64'h84bded03b7cb90a3, 64'h6ecc0146cf66273e, 64'hccbd772e3553ad1b, 64'h5c46b5d6628e538e, 64'h67669f8797feb3f8, 64'h1a0146c7ae648a1f, 64'h4064415a73f3759f, 64'h7c36d84663b1c5d2, 64'h6bfcbe053b46011f, 64'h2059e926944d3561, 64'h9f0210ad32eb81cf, 64'h476d0efe54bb02cf, 64'hd7615d2e34d22ec1, 64'h94836889985a8117, 64'h626bbb046425eb8d, 64'hf62fd7a594cd73c7, 64'haca7ce1485c712a1, 64'hab322cc5a1429bb8, 64'h32d772776052c59e, 64'h7e8110872ead5ce7, 64'h6723399a46c105a3, 64'hdb668f5561f42ae0, 64'h466def9571f6aa58, 64'hb3ef74811fbfd0cd, 64'h3b6000bdb6a237e5, 64'hc48aa554a442d2ad, 64'he301f5a63883156c, 64'hb8d9f901ec2476d5, 64'h342d71d54a80dbd9, 64'h93344cd46296b12c, 64'hb5c0dd791dd0f459, 64'h36955952bbe5ae7b, 64'hf8f2d016ef17933c, 64'he8418e5b2ea88c99, 64'h3305df6b2157f259, 64'h9235ac04e3cbf352, 64'h8fa14b5acb9c964f, 64'h3d3a99c6df258e4b, 64'h3cfb60bf1d24b53a, 64'h7528685e95399dbe, 64'hf8fa639a26055b04, 64'h51bd87142939c741, 64'h6db49c7d555cd749, 64'h8b312c696394e3fa, 64'heec65457cd966483, 64'hdea489db2f1489c3, 64'h9a044fa2438c3d30, 64'he06093ed139acb14, 64'h2960ecb26a40f25d, 64'h7080a64c528866e3, 64'h270e1c542c7ecbcd, 64'h5c4e8693f430b634, 64'h41c70f32c358e727, 64'h4df71c8d18f00a93, 64'h13da3f6c34a6409f, 64'h7ee673ecc56a903e, 64'hbeea63b16492ceaf, 64'h82fe513ad360b101, 64'hd937797e5cc7ae9d, 64'h11060af11b436e57, 64'hc112e2a2516e8701, 64'h838e7d023e1666a7, 64'hdb4e9e1988cf8535, 64'h8e84b8a155239c22, 64'h8ae13b951078a579, 64'h528d01de63b3ff6a, 64'h5425f14524a0e7a6, 64'h8d3a3ccdcd3c2870, 64'hf2393f7687597c1e, 64'h9e803cb055ce6f41, 64'h33cc5c382fa6325a, 64'hbfc43effc045cd57, 64'h3b0b43d973412655, 64'h9e983a3e2e1152a2, 64'hcc7d117ba4cc522c, 64'ha3a73882b84a39a5, 64'hfcec875096f983f0, 64'hdf75bc31747d7604, 64'had1298d2ee100c22, 64'haf656d1658bd46d8, 64'ha4c976a46450ff63, 64'h5d5e3562a272ffb2, 64'h367a426784d13d7f, 64'hf2f3c53e6c23b0e8, 64'h3d59dc9b8085770f, 64'hd9d1608eda3d8140, 64'hd6ac3b2512c10e35, 64'h5016f4e7fff85e4f, 64'h2cb9572f859f1941, 64'hcd9b34ea2d54d299, 64'haefa6b8a8523a99f, 64'h3ea12d30e2df0762, 64'h3b8e95f1a95f685e, 64'hc1cc6745970a9f46, 64'ha6ec06a72c8d3be6, 64'h59edcae19cdef541, 64'h6ee94a6eaf58d8e5, 64'hdc7817e83da73ec4, 64'he8c913236bf65303, 64'hf2598f13a42bf825, 64'hcd9f78058b8bcd65, 64'h8f7987b05e9f5e80, 64'h2f0c2ae96c1e04ad, 64'h439827ad17e33dc8, 64'h51f90bfd3b5697ba, 64'he2209523237f2ca6, 64'h3c228badb8f7a55c, 64'hec9d3d1f4c599b79, 64'h151cbdd5f6856513, 64'hb3bba2db5a8f1db6, 64'h815e9fd29fd247e9, 64'h69ba7c2ee1e087bd, 64'hbe480b39f50ab162, 64'h6441773af0ebf9dc, 64'h82fbf075aa284d8d, 64'hc0cb9ab1d23db98e, 64'h6f1a2cf07b81cd0a, 64'hd4258020bc36b6ee, 64'hf1cdc683fb1a7e44, 64'h3af06f7646b35e61, 64'hbbd63513c35f31fa, 64'ha0c35a11e28d4c2a, 64'h4c7a4b44617a1b03, 64'h86b71a345b9b43ad, 64'h92e7c715b3cb7405, 64'h44e357a8847b2218, 64'hfe50c64e5dcc7871, 64'h187ca2e7d42a171b, 64'h88cb2b361cab0a46, 64'he5ac574471155d0f, 64'hef068b58707faed9, 64'h227093594adf4d64, 64'h64100167c42cbf0d, 64'h3c56ed2e776f0573, 64'he19432d8901a480e, 64'h28c1d37415e2a95f, 64'hb964f446fafd97d2, 64'hcc708dc3c788c70d, 64'hb21b7ed1ceebafc0, 64'h199ab1594f860a1a, 64'hb6e53981e013c353, 64'hb1e7d8a13a4e67c2, 64'hf0b6cab3e8cf965c, 64'h24cd8b1c3e51ec1d, 64'h520bdc1cc138067d, 64'hde3fe5b59acc20a3, 64'h3fea394f739f1f69, 64'h311611bcec2cd25d, 64'hc77cc7ef8a7389b8, 64'h7cdba692277b6ad4, 64'h5c7b69f52cf3add0, 64'hcbc2d9c292c5a7ab, 64'h468bec1d45cf05bf, 64'h4e7edd825a212454, 64'h6d0c9a725769680b, 64'hb317ea07186aec55, 64'h5ebf1907c2debb91, 64'hf2461f63d0a7e34d, 64'h49cc5cc147e6538e, 64'h3dae4aede3cca607, 64'h4915da7bc5f69e15, 64'h4ea6e54017f08c68, 64'hc00706d6be49d6d6, 64'h2559a5d55e68867a, 64'hf39b903d371b9624, 64'h24cd281f9eb47680, 64'hef700470301b56d8, 64'h8b1f79afb428e967, 64'h393d386f12b3ced0, 64'he50b406518749bfa, 64'h4dca3caaac677788, 64'h549680e112546f4b, 64'h9a1bc2be59dec1f1, 64'h345d0623f91ba58d, 64'h3797e56abe895873, 64'he5c61826de1774eb, 64'h3c38c11448d5842d, 64'h1468334def898d4a, 64'he4e8b9a09ee97101, 64'h2a3f8c7c39a675d2, 64'h9a7871f84c65cdf1, 64'h580a8eb439097675, 64'h3d8083e67f389882, 64'h8a5ea82a8ac777eb, 64'hff5035352f1a5df5, 64'hc57b13f5ce806a20, 64'h9c5f2fd77f0ea241, 64'he66c21f2d6c36486, 64'h1c11e008f71db8c8, 64'h11c2f684998d3e1f, 64'h9962263fd840495f, 64'h6c54f48925d98d0e, 64'h9b9adda815f68798, 64'h66d4bb47fc79dd45, 64'he081c6153499665b, 64'hcfb7dffbd2a3a697, 64'heec50d3245da2b58, 64'h87c08fc8d6962a3c, 64'hb028fcde9e8b6fc9, 64'hac7964fa493e6c80, 64'h16212ecdc0b3a55a, 64'h5e6e16fa6a6bf172, 64'ha3072160adb83860, 64'h40b21bc4d63f60b0, 64'h6b3fe4d2a79e6060, 64'hf7f05140978c7760, 64'h66238025a48d8603, 64'h886e2b4f7c91ff26, 64'hbfbeb6c5ede1e754, 64'h83066f8e252cdc49, 64'h98b783b84ac9c7d2, 64'h197faab9cd275595, 64'h5176e166ca7f360a, 64'h852b8eb65c4dfb2d, 64'h5b5db9421a160053, 64'h904186a7d5a701f3, 64'h242287cd2a0dd8cd, 64'h8f057bf2ae6f1ce0, 64'hb6bd319b5b2c5749, 64'h1911110a737ebe4b, 64'h4640276410447ec4, 64'hb4926d1cf47eb8f0, 64'h6de05d3b581255e4, 64'h94e682e9dc796bdb, 64'hcecacc70b45773b4, 64'h77b4a8e2b5b44425, 64'h43d898fc54257c1e, 64'hcaad4c60ef31fac6, 64'h3d9ca43a570e20e6, 64'h117d8f0f77932f32, 64'h4278877ba9f1237e, 64'hba4d29532c81b3e9, 64'h23b6ed70e9853a08, 64'h6d6ad44090044f96, 64'hf72d8fcfc62c474d, 64'h5e213226249a94c1, 64'h90a550cb60ab8c17, 64'h153459ecc9139970, 64'h6c60d123991df8b2, 64'hc560d750f1cdaa5d, 64'ha2f515a25bb1f0f5, 64'h2a6b19c421bd9394, 64'h5cb9cd18ae99f4eb, 64'hb6d6249341da3247, 64'h23defb8359529336, 64'h936afb21c51ee7a1, 64'h8f1e255254e04822, 64'ha5cd9a2a4f8f9069, 64'haca573e2da0e36af, 64'ha958f43f97c065c0, 64'h59b6cfabe26d2e6c, 64'hfd513773ca985615, 64'h99acadba31e833c4, 64'h5b953d39680bd628, 64'h560e0ada7b075748, 64'ha28d4308431978f2, 64'h4bf13d432aea8694, 64'h59d23e30876338e5, 64'h858dca51fef0438f, 64'hfb774f6478c66aad, 64'hf948f26f43749b74, 64'h91de779e7cd310d4, 64'hf839e403d8aeaacb, 64'h43652fe4797d484e, 64'h386f39a38efb1e44, 64'hce6fb2ca189c6a38, 64'h3ded16e6fa96deb1, 64'hf69762f19594fdd6, 64'hab0fd05e514d6512, 64'hf48079f0b0bef6d0, 64'hb008aee812aa3056, 64'hdcb677b3cacc5ce6, 64'hb461bafac1c9a275, 64'h3593cf4dbc818a0d, 64'h273c85eeb9aaf95e, 64'h10a1b293ca4a1566, 64'h85f94600410d8771, 64'hbf04e9795bc1ca35, 64'he41dc0b33b418c3c, 64'hf1408d5df8fae39c, 64'h591392cadeff2a16, 64'hda1f7c2e75e83475, 64'h6748c52053c8f557, 64'hfe6077d24d6157d6, 64'hecf64f0976ccea61, 64'hf080a2bad952a06a, 64'h3562f57a99d3f824, 64'hb1a4067571659b13, 64'h112ba5475e145b5e, 64'hd958c7121f13e7c5, 64'h294cfd3eb86dd088, 64'h8b65e24c878f5ea7, 64'h69aa94c5a0d7e06a, 64'hdc5a3db552762711, 64'hdabe235d73fd149b, 64'h883c752ebf1c0f76, 64'h4e17dc99ed315f4e, 64'hb87f25dca48b15d0, 64'h5185a9b9b700edde, 64'h4dbb462fd3f2da21, 64'h12c0de1e37f812a5, 64'h95e10359baf28b6c, 64'h863202eae2ac9da4, 64'hfa3572f07f6d2edc, 64'hc8511eba86beccc7, 64'haf9fab4045f8519b, 64'h2a4a3e3dfaf64f23, 64'hd399459b547df6d9, 64'h9c994bc36b37932a, 64'h3a52359074853b30, 64'h575337d413fd6297, 64'h6cf7e8a6ed04e51c, 64'hd6c49fb899c72729, 64'h5c79a9d34780e0d7, 64'hf571d7de9781a4fe, 64'h4439ab7c4be02d5f, 64'hf64d97384950bd88, 64'h299c837b3c269f20, 64'hc7e4da26ba1a79d4, 64'h791b26e1ce835953, 64'h8c33fad573437895, 64'h2c2fa1f0e4237ef3, 64'h52247275a3e70f11, 64'hfc4c94e63d75d7e1, 64'hf7a52675aca6d50e, 64'h2ee54511c9433430, 64'hf46d1a9497113cab, 64'hb540d4dc1652d04e, 64'hfd60cf645c6e0165, 64'h15bca5f1d20e2e71, 64'hf994a305c1057024, 64'h10a816831f34dead, 64'h9c39832460925613, 64'he3a3d95ce1ae3efe, 64'hfd012969bbccb758, 64'he273bc0a5cb74d8a, 64'h2aaeb641dfaff87e, 64'h58d55b3f74a3c6c3, 64'hab0c1958a1394a73, 64'h750583aa6cad1664, 64'h2d7185f290207964, 64'h47e28e45c52764f6, 64'hb1f80c7821433156, 64'hfd6c6c18cb4f462d, 64'h46ad9f5c1760d6b9, 64'h82cf2a5264a87ed0, 64'h9329aaa2ae51c0e1, 64'hcf552f5a13402a28, 64'hbb6e50fe56e01710, 64'hfcbc9302db191789, 64'h967f0c6f9f76b946, 64'h3e19211e464ce5ca, 64'h34f691d76aacdd47, 64'h2ade8ae28ab49b4a, 64'ha93c15e92d54ba81, 64'h629b6c9f20e22c7a, 64'h8e2ec471ac11cdad, 64'ha3b69bbed354255d, 64'h48893088a45d17a6, 64'h58adc8c3254de34b, 64'h594343cb2120244f, 64'hf60eccaebe850b59, 64'h2859c14fccb4631e, 64'h64846ce3eabe9335, 64'h86eb5cc6e1723dac, 64'h44ed59c168204be8, 64'h680a7634274fd4fc, 64'h5f7186dfae549203, 64'h7ff86e9fe303fcd7, 64'h50b88a8a652819ce, 64'h5ce2914e946ac7eb, 64'h3d2c336e399420c8, 64'hf179c4f96a653c4c, 64'h9ce74f361d3c8b4b, 64'h31ce50ba272044fa, 64'hd2e8616928c1569d, 64'h8bea75363556b4c0, 64'h52ea8060e3d3112a, 64'ha7951ef6f7476fda, 64'h9fee735d1248e431, 64'h73c0fbbf1562d247, 64'h5b5b327783970927, 64'h9a1c38d04946ab21, 64'h95fd209c6ec7e49f, 64'h899468dc3f0836a0, 64'h359ed1a5c5158663, 64'h5f318e21aa9b6224, 64'h97b59784e7e32df2, 64'he35d33957a58c3b3, 64'h4122ec79a7b9e649, 64'ha8d733ccb62e21a4, 64'he9cb2751cbd1c67a, 64'ha611e007a03b5381, 64'h430fea49ac53e34a, 64'hd37ae3f8ed5b7e44, 64'hebfefb9f96a9e920, 64'h4e5c3311601c8409, 64'hff76850e8e24ba66, 64'hd3d14e559f48acb2, 64'h89a9cd9263a64623, 64'h91109f0b119dc7c9, 64'he267937296c1babc, 64'h15d3d9cdd45ca807, 64'h307c2c7d175a710e, 64'h7ef5e322f68ebf53, 64'h2677a8d11fbe5f72, 64'he32f3de7d5211926, 64'hd4caebdb8046bda9, 64'h76991d437041a2fe, 64'h9bbb4acdbef3f53b, 64'hcc3ae690ad26dcb2, 64'h96fdebd172f966e0, 64'h5cc794d854b3107c, 64'h571518fbb3dc560b, 64'hc6fc62e19f6dc27d, 64'h457cc1ef3ea7a14c, 64'hc7c3c151fae2f2c0, 64'h13d1820f4bbc4d46, 64'hce27b3eebc998412, 64'h4b090234952c9681, 64'h9c8a6425bd21d997, 64'h7f481ce27129e3dd, 64'h59ec1a164931b308, 64'h26336805ab031349, 64'hb0b2688bb4f6620f, 64'h10c145e8792e442e, 64'h2d69adc28e62e0aa, 64'hfb2333cb87d3945e, 64'h69ea7ea7d3525443, 64'hf85e4bdf54e8dc3e, 64'hd0b8528cff12ee0f, 64'h2ad67b368f738caa, 64'hd33f12b36a4f83c0, 64'h7afc630cc437740a, 64'h279a66cb6686bc77, 64'h974a1cc24942b2f3, 64'hd996c27ec7cde28e, 64'hf7baefa48d846328, 64'h2990e000f0c9bffa, 64'hd837758e92a90d44, 64'hd8b66974e39b1710, 64'hca426cd39919d828, 64'ha3abf416daa75d12, 64'ha554fd7a418e20f2, 64'hb5f50c7b8faeecc1, 64'h4f2de6391030533b, 64'h4884fb83b1a7f01c, 64'he2cbfe3ad75e5da9, 64'h29f21e272111eb33, 64'hc6c83b4d545c2992, 64'h513b945e107ae603, 64'h27a63ca0308b1525, 64'h363f17517ae01158, 64'hd3648125d2f398a2, 64'hea65c32a7a764b7c, 64'hba172c7285333f8c, 64'h1bf653a8234db512, 64'h4b06b274fb96d6ca, 64'hb60f6503505262c6, 64'hb980d052aeb91b44, 64'h1a63bf5c66c1cc16, 64'hc9b1d8e922d872a9, 64'he4408f65ef688c52, 64'hdcbd92ea2c2bae15, 64'h97a4423cb9d07bb3, 64'he51d7f2a26fc7ab0, 64'hd3c8f1d952b952cc, 64'h9e262312bcc03f97, 64'hca7c0e7a56b83555, 64'ha1c536ed54fe555a, 64'hff9894c6d37b397d, 64'h735acd9de2fe7ef3, 64'hbfccde57eee63620, 64'h392fc2d556c2a9a7, 64'h267f2e6f5c50c12d, 64'h6b7c3a7ba7d9dbc3, 64'h812a2f5dbc3d950a, 64'h509d180a39889ad6, 64'h6afd4af07923b939, 64'h754f74d2eb41b8b8, 64'h50b23297647d8bf3, 64'h43a67b456942f328, 64'h6d90b7199a1a3d08, 64'h52cebe8a4e47351b, 64'hbc9321d3ea71613b, 64'h2d4da0ec3bbfd599, 64'h2ff241b0b410db25, 64'h435cc2aca118e11b, 64'h40672438d4430082, 64'h5bdd9f49b0b54108, 64'h33b230ab596d49cc, 64'h575683b0a86b4fa2, 64'hb3694cb2dadc13ac, 64'h3c00d57ec680ce03, 64'hbadd8e9095cf7f83, 64'hac0a038e25994c94, 64'h33400cd573bcb9fe, 64'hbaba9d773846eeab, 64'h6d5ae0da8781cca6, 64'hf06935a01d3f41ed, 64'hd6f63862fc32c7ec, 64'h50253ab9e59d1eea, 64'h55ac0a60cfc3054c, 64'h7e5da2ff9f6d134d, 64'h48ccd7f9b5071033, 64'h33af32bc96532375, 64'h86a391cbd8edefb8, 64'h838d6cf4cc55dec5, 64'h7012150c59e5bd95, 64'hccef3c3a746e71c3, 64'h87394e8b9a8eb243, 64'hd4b843509b844c9c, 64'h71796b82368a746b, 64'hb881b7f5e3f9d317, 64'h2a02cc837fe42fca, 64'hf049dc88973e00d5, 64'h92dc603c1f3bf013, 64'h9078d7d2ad170489, 64'h332e9a5ef5870c83, 64'h3f138132b1be0357, 64'h51d7853e2a05fd8d, 64'h4e9dbed2603249e6, 64'h7f892065483edc22, 64'hbe99d6bcd1b9d242, 64'hcdd58a67bbc79740, 64'h50b6e18d428286d5, 64'h2a30d8316f34163e, 64'h24f1a992ad4b23f8, 64'hf3f57d0fc55a1bd8, 64'h2c0dd3e514ea5e31, 64'h605f91d8fe4a4fa3, 64'h5b1461f2c1007aab, 64'hbbf7909e9969f056, 64'h683c2c7e41fbd821, 64'hfb3326e11fd08363, 64'h48b1d5455a22c892, 64'hea47e2d4bb356854, 64'h4fb0724d377af5c7, 64'he351c2d7ce820921, 64'h1936861ae3083e6c, 64'h9d1b04997dcf15dc, 64'hb1b9759619775d95, 64'h5f46ef4c2521b1de, 64'hb412af936f85d6fd, 64'h82f2f07d558d8465, 64'hcd30d0b91b29bd3d, 64'h53785c179dbe35b2, 64'hcda1cd6aa0624361, 64'hbf51394c15a58e1b, 64'h4d2e815e1a1a1e24, 64'h8800c303fd64c7a1, 64'h133f507e79cf9bae, 64'h112613d9a317e075, 64'h3c018f65bb0edaef, 64'h3650cdf9d6dbb032, 64'h417b961d64882afa, 64'h4756bdc7d1d8229e, 64'h85aa2fa3e1b854a3, 64'h2f387b7087bffc7f, 64'hca632445fb7d8d83, 64'hb19c53e73beb97ae, 64'hc658734d21e9966f, 64'hc710bd7cd6acf7c1, 64'h9635d8508640c48e, 64'hf0c43eaf1005f4e8, 64'h124bca3d4c77e53c, 64'h895cc30d91b332f3, 64'h691c34e056402fd9, 64'h40917324d01151d1, 64'h5bd24da386313ba8, 64'hd2b5b65fa2f7555c, 64'h7210e7f03a74fed4, 64'h6f6fbe9284737728, 64'hfdbd84735434f20a, 64'h37c0e6d844f028d9, 64'h42c08dbc22405ec0, 64'h6793edd354560ef9, 64'he5057495cb432683, 64'h2a2cf372dc1eef4d, 64'h2a4dbd09bcd99060, 64'h997a532b24d581d4, 64'he9475ac3e1e55ddf, 64'hda86401968b237e3, 64'h45822281ff4e8a43, 64'hd42944e91a1c5aad, 64'h6996315dd2ecc48e, 64'h8ecff4ae4b4fb7ca, 64'hce4b08d24ed1fbf1, 64'h101879fa47843c01, 64'hfe68abaaad7cfab1, 64'h44f5d974b4ac6c5d, 64'hb4dd672da9c73c5d, 64'h20ee80394a4fb722, 64'he1003cb5c05679d8, 64'h38469d8c57a95625, 64'h970da436d658d3ef, 64'h401fb8cd286650ce, 64'h6ba6064beaf6ff46, 64'h4e85f35d29fe382d, 64'h1d6d22c36466a393, 64'h1907ccae9bed9aa8, 64'hb169e3f37e841c9d, 64'hc1de3831883ef94c, 64'hb8908b87475a93c8, 64'hc2b4fc88886496f7, 64'hb949dc657b351cbc, 64'h896cfdb619f7ebf1, 64'h856f29af322624e7, 64'h3232f1e178010c7a, 64'h9a4aa2fe6254e96e, 64'h36849a73c1f0418b, 64'hf72458a3c012fb68, 64'h227ed38ed9d165b2, 64'h2034103278b70324, 64'heeed54954f29c91b, 64'h2eb57161c6eff33e, 64'heeddaed85e2f3637, 64'h47ca39bd3bcbe85e, 64'hf72d30c69a646e95, 64'hde6bcaef5a00b749, 64'h1d8b744c7ce9baa9, 64'h41b4d8248c8e5b39, 64'h911df5d956a1116d, 64'h59c9f76e15cd3afd, 64'h74e57fef5daf7a43, 64'ha4ad792ade57d7c3, 64'h863bd42523d9990c, 64'hf0090a14d1ff9bde, 64'h67b979fc5f5ffbfb, 64'hf11aab7869f9821f, 64'ha897b036fc7b8e5f, 64'h18d14a885b82ed64, 64'h477f1f6ded5e21a1, 64'h9445d73a1ce428e9, 64'hc54273d4b42e1c28, 64'haeebfa18f55ff9d7, 64'he1e785b1c4c7c571, 64'h457098a3311fa3a8, 64'h45036120415286a0, 64'h984fbde0af21699a, 64'h8e94884f1d861b4c, 64'h6728b5b8f8412c0a, 64'hb6ec3b3068bccfe3, 64'hb130b5e84fa056f0, 64'h229838b78ebc71ee, 64'h558b6a448398b146, 64'he87a8c43ac6aed9b, 64'hbd98ba4b289eea87, 64'h831e315b710ac408, 64'hab3ee8b4550e7259, 64'h6bef7ef5fb71abf5, 64'h2b8df6173ffa56d0, 64'h495eff10b7326f20, 64'hbb48ff10cc5757e3, 64'h6b735dccdc93a873, 64'hb75cf8aebb2eb028, 64'hd546fb79a6f11e14, 64'h7555aa481764476a, 64'h9ee8cbc4974da23b, 64'ha031a5155d7c1dfc, 64'h952bf2dc39329037, 64'habf75cf821339e44, 64'he204bd3643df8403, 64'h5685cf78e4563c7d, 64'he40fe5e5d8b441fd, 64'h5e76eca0e8900dfd, 64'hc93b8877adf09e4d, 64'he7f3e69fcbf39900, 64'h75f09c1f5dd23db1, 64'h6e87df6f1ebd29aa, 64'h673931af64bb010a, 64'hdfbff7f1e549bb26, 64'hf721eb945ec48fd1, 64'hb6659723a7ef976d, 64'h4a2fbe66e0cc0a2e, 64'h43626bf5c3738c5f, 64'h32b826f729a2ffeb, 64'hbce098bb8e50fc2d, 64'h7a4cbfaacac36a02, 64'h6619310ddccdcca2, 64'hf6ebe0d4fafd7868, 64'h52a176e7739a0846, 64'hbe009b78e6c49020, 64'hbab6f461c5f3a5c0, 64'he404520568114cbd, 64'h9235f6139058446e, 64'hab6b7947e6d818fb, 64'ha032d713f8c90615, 64'hbfb6689373ab825e, 64'h9b7925a2ed5b638e, 64'ha470a9e1ba62036e, 64'haeb5c84f60acd654, 64'h40cce4bd71e00747, 64'h342f4c01d651eee5, 64'hba82b33a7040e46d, 64'h3921c0bbe2311c88, 64'ha960161eff2f46fb, 64'h284374504ac37bb3, 64'h2413c258c2bcef49, 64'h364c4e99e399296a, 64'h85f4808b8e47d6ea, 64'h1a347251a35f7494, 64'h46a0a714433db0f6, 64'he6e05f75e51f8a49, 64'h11437e31d7c0c15a, 64'he88d3da18ade106a, 64'had7b51c3c844c09f, 64'hb4816e9b7e301ce2, 64'h99a0e7b799c63624, 64'hda1c7fc949b4bd10, 64'hc5bbfe7dd2f5fdf6, 64'hcf49ab14d1d99183, 64'hd706f6ef74342af3, 64'ha44af607c54248d6, 64'hc8be6587f610ab05, 64'hfa049ffc97894b18, 64'h7fc70226d886ad14, 64'h44ca6630c7ef7fa6, 64'h3e1531529dfd9900, 64'ha1a3b9867a0ae21d, 64'hdf7dfdfb926f8ba7, 64'h8641503e7459a39a, 64'h1eef1d8366ea767c, 64'h2646935c97c0d455, 64'ha9b86b96c8448acf, 64'ha7cef7563ce50347, 64'hc40efd0493b9ebec, 64'h288558cd15f55f68, 64'h57b2f750b59a85fe, 64'hefde842af7f59688, 64'hc77dd5a956613ae0, 64'ha54bed5447768bcc, 64'hc42a6a9c37cedecc, 64'hc58d8a5ee0761bad, 64'h8cae786a1fc09abf, 64'h7bbbecffd914309d, 64'h3b2400c719411198, 64'hbfd8b177972138d9, 64'h1a183474fc5f59c3, 64'h98a3c82a9c7006a8, 64'hcd93dd35e8a1dfca, 64'h1e94867763a4a6cf, 64'h4005a4e27fa2e8fd, 64'h25f3ca55205730a2, 64'h5836a593e90af8ff, 64'hfa214c94c74af571, 64'h102d858ec073a4c7, 64'h154738463874acef, 64'h1285fb0e33ca5ce1, 64'hb50056e8b87beab5, 64'h690efef1bf7c5d3f, 64'hdb5a5ed22f492a6b, 64'h24fa4e366942dab3, 64'h70ee9c5752564678, 64'hc50017e65d3a8b4f, 64'hd008ddd5eab6c909, 64'h8b27e002770fb084, 64'h25fb95ac51aebbca, 64'he4cba4494b06d202, 64'ha515e03d86cd4121, 64'h26a63fa5e7d933dc, 64'h2043d707b35e59d4, 64'hf94790d4ba3fecfc, 64'h5e37d4f021a029f1, 64'h9b230b4fc00b491e, 64'h661f8015ace67d90, 64'h97fb604a182f7f90, 64'hecf7779b6b338e7b, 64'h6b0e7498db201ae2, 64'h843a08c87c41aaaf, 64'ha990cbee42d33a66, 64'h8ecacb69b074d9a3, 64'h914e70c2ba1a48c8, 64'h9fa61503d9eff4bc, 64'he300406e277b3d9b, 64'h4e1003d91d1e12ff, 64'h46ef1dcabd051f5c, 64'h22d9d1cc353a8afb, 64'hc8fc018c7aa356c3, 64'h55a104a4aa8e6b75, 64'he4dd7edf19067a70, 64'hb657b76fb073c1a9, 64'he052a9d13f211920, 64'hbb11faab28efaf21, 64'h1d971f95b3641bbd, 64'h156ead461aa1bc6c, 64'h18de64cb7fb2d259, 64'hc5e37fa8fe20b866, 64'h4662c6e2ce2bd74f, 64'hcedbe7e9e1569792, 64'h5b6be3572fe6ea57, 64'hcf3558579830f28e, 64'h738456571e12f1d5, 64'h1192dabc5bd87b4a, 64'h51266d83822c75ad, 64'hedaab68674011847, 64'h551795c5dadbf26f, 64'h59aafff7ebbd7b7b, 64'hdf38060fa9510d0a, 64'hc37129f535c1e99e, 64'ha0b0985d5e7d2bb5, 64'h8548612f4617aebc, 64'he878479c72c4a2a2, 64'h826a8a4dbd22fc33, 64'h2d53c5ae88bc510c, 64'hd327caddb28fe246, 64'h5d32387aba8f4830, 64'hf043f80de6bf0d56, 64'hc222e7c84fdd417e, 64'h6965a05596053274, 64'h6b73a4ec7d611654, 64'hce723be828f214ec, 64'hf984e8e7b91bcba2};
    //parameter [31:0] RANDOM_32 [256*9-1:0] = {32'h7415d4fc, 32'h100706f6, 32'h3338ae94, 32'h3cb3d3d0, 32'h6f3964c5, 32'h749b4f9c, 32'h41118bd6, 32'h1692b199, 32'h74273502, 32'h31b15f9f, 32'hd02dbf0e, 32'h5b38c811, 32'he255597a, 32'h24691dc9, 32'h38c26188, 32'h279a6df2, 32'hf5e4bb95, 32'hb60cee0d, 32'hb4c29df4, 32'h1463a1bc, 32'hfd53a014, 32'h534e7a98, 32'h28c634b3, 32'hea101b93, 32'h5510eab4, 32'h14a5e7e9, 32'h42ca6e74, 32'h85fa4142, 32'h99c9c923, 32'h9d6eeea4, 32'h288f6d65, 32'hb6a7f219, 32'h1bfd23f9, 32'haf4f8b03, 32'hf2b3e6dd, 32'he8d10381, 32'h316d2387, 32'h6f7143cf, 32'hee9a208f, 32'hc431e548, 32'he3fe5385, 32'hc439e735, 32'h50c85ea3, 32'h76bdec37, 32'haf39d87b, 32'h2b89fe1a, 32'h7bfa99fb, 32'h71f3ecd8, 32'he8cfa344, 32'h10b05a58, 32'h5e651012, 32'he4a04858, 32'hea0c6651, 32'h13cc0ea3, 32'hb5d0b4e5, 32'h395c99d1, 32'hefd2aa4e, 32'h1fd70cf5, 32'hc4ee272d, 32'hbac414c8, 32'h14c56f78, 32'h16cb2690, 32'hde681dff, 32'h94ad61e4, 32'h2dcd3560, 32'h9c950cb6, 32'h96a5b25a, 32'hd026df15, 32'hd1b48b11, 32'hdf4002f5, 32'h957f6665, 32'h1e6157c5, 32'h1ab14476, 32'h462b94ef, 32'h965502ea, 32'h21461989, 32'h985817a7, 32'h4c8ee4cd, 32'h3ee72ff5, 32'hf8ce0734, 32'h49903f0f, 32'ha4ca1450, 32'h35a14367, 32'h20ce2918, 32'ha184e1d3, 32'h5c2abf16, 32'h9b238bd9, 32'h943a4233, 32'hb09dab42, 32'h1feb9cbb, 32'ha721d7f9, 32'hc4a94d1d, 32'h4e79c279, 32'h3e6c9a32, 32'h8debbe6a, 32'h4f30f41e, 32'hc06a73ea, 32'he9e034bb, 32'h13592f45, 32'ha406dcbd, 32'hf40ad21e, 32'hebbedaa9, 32'h6d9a12ef, 32'ha108d609, 32'hee48963d, 32'h6ec5285d, 32'h39bfd60f, 32'h306b4373, 32'h152a7bea, 32'hd681f97d, 32'h3a497f7a, 32'h2f707237, 32'h62bc9eb5, 32'h9baef383, 32'hdabc7bfd, 32'h7e5f0b25, 32'hcfaa3464, 32'h85a92d2b, 32'h13ba5d4d, 32'h7815132c, 32'h5ba8a406, 32'h9aaf8c1d, 32'hcd1a5f44, 32'h1cf02f89, 32'hb2f9fd44, 32'h1018b34f, 32'h6a611834, 32'ha121c1db, 32'h99ee465d, 32'h5489ce87, 32'hc4015651, 32'hc5383fea, 32'hdf799dbf, 32'hb0fd4369, 32'h6bb464a2, 32'h705ae7d6, 32'ha542b9d9, 32'hf9b66651, 32'h3fa8224b, 32'h62673167, 32'he3331849, 32'haf0d815a, 32'h4c9168ff, 32'h8ea6c9b2, 32'h9965b1cb, 32'h8c90130c, 32'h9886a28d, 32'h623ece78, 32'h6ab3a95e, 32'hfbe04892, 32'hd2d89930, 32'hb5381c38, 32'h36a215c8, 32'h62d75eef, 32'h9e33ede2, 32'hebe9d02f, 32'h4db55915, 32'h3e4fa159, 32'hbedc4daf, 32'h4b872e8d, 32'h73cdbec9, 32'h48147296, 32'h8bce4150, 32'h34a42555, 32'h928ffb51, 32'h32b0e0c4, 32'h454ab2fc, 32'hcc789686, 32'h5dd8d45c, 32'hdabaf553, 32'hdffc6991, 32'hd6567229, 32'h27b2cb6c, 32'hb8d81571, 32'hcfe85c98, 32'hc8db77c6, 32'h4e53de8a, 32'ha7c0b741, 32'hcf2e688c, 32'hcbdc1fc2, 32'h580f420c, 32'he85063ed, 32'hf9f00c63, 32'hfe8a0428, 32'h8e579c01, 32'h655e8695, 32'h367eae0a, 32'h174bc1c8, 32'hdef68dc5, 32'hb5d37c37, 32'h7a0e9959, 32'hfd8a584d, 32'h4b74b5a1, 32'hc40a97d4, 32'h1da9bea5, 32'h42ded520, 32'h575c0a43, 32'h9e6c7d5d, 32'h6b71a174, 32'h8aac884e, 32'hf643a50b, 32'h17c1ede1, 32'h7f99b0e8, 32'h4524d3c4, 32'h238dc2aa, 32'h2a2a1ce5, 32'hd0b60fb2, 32'hc7e406fb, 32'hdb011d79, 32'hd5c32a9c, 32'h326be981, 32'h14665b8b, 32'h7e0f63b8, 32'h16ab024b, 32'h6ec39d10, 32'h7c93c0a8, 32'h82bcc65b, 32'hd0c25b12, 32'he91feaee, 32'hc9bad6f2, 32'ha471793b, 32'h914542a0, 32'hf44958a0, 32'hcf08357c, 32'h32ef1905, 32'h3d08170a, 32'he964ef79, 32'hbaab5d27, 32'hea3af978, 32'h4bf6d368, 32'h2cab70f1, 32'h333aec66, 32'hd494d6d2, 32'hfbc7ba64, 32'h9013a95a, 32'hea95e1fc, 32'h780fe9a0, 32'hf1552f68, 32'hbc0d066d, 32'h168c86eb, 32'h5e3cd065, 32'h960b41c4, 32'h7caf51ad, 32'h559f8cf3, 32'h9a6be279, 32'h8c24ebd8, 32'h765a9c6b, 32'h691c49e8, 32'hf0d93180, 32'hecd97cfe, 32'h24fee82f, 32'h5b734c9f, 32'ha1b3dd86, 32'hd3eca30c, 32'hb8734b43, 32'h99d00555, 32'h1dabe489, 32'haf627605, 32'h8c905792, 32'h98f8c82c, 32'hd40a595e, 32'hfa3cc4b4, 32'h9ef226c5, 32'h26756074, 32'h7c6a7c13, 32'hfa158191, 32'hf97811d5, 32'hd5d12c41, 32'hb07ef100, 32'h13271908, 32'h8618e439, 32'h80788680, 32'h3109ffb2, 32'hc5fc9dc8, 32'hfc4084e9, 32'h614a389a, 32'hc52c87f8, 32'h2df518d9, 32'h8915a865, 32'hc8d60369, 32'h157fe7da, 32'hd265b4d6, 32'hb1648c19, 32'h7bd1b876, 32'haaa58b89, 32'h844348a1, 32'hd74bbfe5, 32'hb1b007fb, 32'h51c9eb43, 32'hb13713f7, 32'hdd66184b, 32'hc35b63fe, 32'hc9b63a6c, 32'hd1d8fd82, 32'h43495002, 32'h5a12f616, 32'hc2ac6e37, 32'h43630cb9, 32'h323453a1, 32'h1664046a, 32'hb1e536b0, 32'h2353bbf2, 32'h41d4854b, 32'hbab729fc, 32'h591595cf, 32'h787932b3, 32'hb973d2a7, 32'h2e4a594a, 32'h365c2df3, 32'h777bce9a, 32'h33386936, 32'h3d4c7f36, 32'hc5088ec0, 32'ha03aa107, 32'ha92c2858, 32'h56ea6e80, 32'hf2dfc025, 32'hcbb94037, 32'hd8771657, 32'h6ed2c06b, 32'h23399161, 32'h68d645ce, 32'h869680de, 32'h418c8992, 32'h89e6b592, 32'h65b1dd82, 32'hcd032f5f, 32'hfc91f33c, 32'h996091f3, 32'hcce86cc3, 32'h8eb26ba2, 32'h33fbca5a, 32'h43fcf617, 32'hbd7fe8d5, 32'hdedf39ae, 32'hde74f60d, 32'h70c5dda6, 32'hbc101e2d, 32'h52bd8b9f, 32'hf022f9ec, 32'hbeec9911, 32'hb9ab6447, 32'h69f860c3, 32'hc4265bb2, 32'h7072a473, 32'h10bf4106, 32'he723d608, 32'h2cfbef91, 32'h5880d2bc, 32'h925c253e, 32'h3134831c, 32'ha3543d61, 32'h7dc435a6, 32'hd6c0a2f6, 32'h62f7bc4f, 32'h4527db86, 32'h5b8b342f, 32'he291070f, 32'hcc451056, 32'had7ebaeb, 32'h77ea6240, 32'ha150a13d, 32'h8920ce2d, 32'hda4bc425, 32'h9995d92f, 32'h8c495245, 32'hdb816573, 32'hb82c9b92, 32'hf3b88066, 32'hd91d5db2, 32'hfd710d95, 32'h5d4fa328, 32'h122537ed, 32'hdeb0d7d3, 32'h4d60fc16, 32'h82afd770, 32'heeaf0ac9, 32'h85f888b6, 32'h74756f15, 32'h6f848b7e, 32'h3d7e0e7f, 32'h569c9ca5, 32'h32a2bcfb, 32'hbbd3b42b, 32'hceb2e4d7, 32'hce097c14, 32'hcaaf02ab, 32'hab770718, 32'h5d3c9e5a, 32'h7212abce, 32'h71a9498e, 32'h5ce06b5d, 32'ha8b6a5fc, 32'hddcbd8fe, 32'h4c7ce996, 32'h77e7bdf3, 32'h5f443709, 32'h5079dd16, 32'h56de8b25, 32'h8519e57f, 32'he5367669, 32'h9c7bcf30, 32'h7b117123, 32'h52f53348, 32'hb3c9f4b8, 32'h134de040, 32'hf13c53d3, 32'hcb237d51, 32'h62119510, 32'hbc06661a, 32'hb53d4675, 32'hb62a9b1b, 32'h75ea7113, 32'h65461e3c, 32'ha7985e67, 32'ha342e3b0, 32'h38c92851, 32'h8b66ea29, 32'h3c261976, 32'h76f19a45, 32'h36c338c4, 32'h4ed9ee9a, 32'hd01469c7, 32'ha1af07a9, 32'h8a4ea40c, 32'hde50f460, 32'ha808a4b2, 32'h80f0eb59, 32'hf3978053, 32'h3469f9e1, 32'h97c247bb, 32'h76ba9f44, 32'hdbfe2664, 32'h9b0be95f, 32'h1f899fe5, 32'h1cb7fc16, 32'h7575ec6d, 32'ha5ae4f60, 32'h544f4a90, 32'hb8d83a4b, 32'h6adbfddd, 32'hc347fa09, 32'hcedf4dc1, 32'h8e292173, 32'haa9d9d85, 32'h47025b5d, 32'h6bcaccf3, 32'hfb137511, 32'hc9dbc234, 32'he56436d1, 32'h4aecaaf0, 32'h1a72bec4, 32'h9589a412, 32'hfed003c3, 32'h8c027052, 32'h99150995, 32'ha76e221e, 32'he1fa0344, 32'hba07d5fb, 32'h86c328bb, 32'h34303186, 32'h322212e4, 32'h827badab, 32'he4a3b722, 32'h722e8a6d, 32'h21486b61, 32'h162e4b41, 32'h88d79fd2, 32'h2a407c7b, 32'h87fbd84b, 32'h327736c6, 32'h6fcffdba, 32'h3e008eb2, 32'h55abe8b1, 32'h1403017c, 32'h6b75a597, 32'h210539fe, 32'h13fa6c19, 32'hac6deee1, 32'h5d0bdb54, 32'hfe6e35fb, 32'hb7e8d92c, 32'h1988ee87, 32'h81c2f24b, 32'hf0f0c447, 32'h91840a95, 32'h7b3141d9, 32'h4cdc100c, 32'h5ece8619, 32'h44d4b4ab, 32'h32453824, 32'he0d894b6, 32'h6ca41621, 32'h8e3145e6, 32'he1ca4c28, 32'hd30072e3, 32'h8eaee83c, 32'h951ec274, 32'h5acf06fb, 32'h5e3b6cdc, 32'h5e31c3ad, 32'hc468ec21, 32'h80accaa1, 32'h19f43a99, 32'h18e833be, 32'hb0e24e54, 32'hc844f46d, 32'h1990fe70, 32'h3e6b80ea, 32'h1c8e1b81, 32'h8ae50790, 32'h77c3ed81, 32'h7cf9636f, 32'he1894e9b, 32'hd5854e8c, 32'h1c380e8e, 32'h1f33d238, 32'hdf51a9a7, 32'h818bff97, 32'hc97e1766, 32'h1a63cb95, 32'h49756a21, 32'hf288c358, 32'hf9a310d2, 32'he77bf2b7, 32'h48987389, 32'hb4365b68, 32'he0e6e739, 32'ha12eb503, 32'h4cd34b77, 32'hd38233d7, 32'h2f52935e, 32'ha4672b93, 32'h4b96fb7e, 32'he171d686, 32'h1f76984c, 32'h40cfb7e8, 32'he39ffcb2, 32'h9fa1abb6, 32'ha5f50534, 32'h53b6a5d1, 32'h983ee4d6, 32'h467af39c, 32'h497793a9, 32'h36d7ec6f, 32'ha08629e8, 32'h62f687e7, 32'h9fc1a7fa, 32'h1e33d8fd, 32'hf391fdd8, 32'h3e36a456, 32'h11c1ad70, 32'hec39bbe8, 32'hdd3ee41c, 32'hd56b33a3, 32'h5d096722, 32'hbd1ce0a2, 32'h2e6aa459, 32'h18a8098a, 32'hcd3139a0, 32'h58cd8ede, 32'hff657a5c, 32'h566909df, 32'h89b56ada, 32'h9d16d34a, 32'h5944e9c2, 32'h4aaae295, 32'hb700c957, 32'hf90f5bf2, 32'hd17aaa2c, 32'h2336f24b, 32'h7af6257e, 32'h7bb26acd, 32'hb3984a20, 32'ha476d463, 32'hc697b3f3, 32'he8fc1664, 32'h3a6726b5, 32'h5cef7e0b, 32'ha33f0802, 32'h76a3be65, 32'h2b9bc04b, 32'h3e8601c0, 32'h9fe9a2e9, 32'h85ddcbc9, 32'h486b2b85, 32'h3fa97643, 32'hbf0e31d1, 32'h5f4b44d7, 32'h76d38178, 32'hadb21986, 32'h402cb266, 32'he6a9ed84, 32'he106e5f3, 32'h5f29a662, 32'he7d02299, 32'he2dc7036, 32'hdbf1cd45, 32'h62a4333f, 32'ha87d311f, 32'hd53e6cf4, 32'hf5832a2e, 32'h3f7ad8a7, 32'h60d1ac96, 32'h6b41baf7, 32'h8c83554b, 32'h21e5d4b9, 32'h2d9edad1, 32'h73573c3f, 32'hef307939, 32'h6ec590f4, 32'h96a0b108, 32'h84ed319c, 32'h4ee1430a, 32'h15585c97, 32'h3d3b7f9d, 32'h6540109d, 32'h2d771ea1, 32'he5775880, 32'h5a38190f, 32'h469f9ae5, 32'h40d2f964, 32'he18aeb2a, 32'h80eb6092, 32'h86ff92e7, 32'h52250dfd, 32'h6ce09e5a, 32'h4d10ad51, 32'h6bfbb4f0, 32'hbc3908d4, 32'h2c5dc152, 32'hc297b605, 32'h4a4b4225, 32'ha9348d09, 32'h20328b95, 32'h7e63bdd7, 32'h4ceeeab9, 32'h76e92cb6, 32'h2e694533, 32'h230abf33, 32'hc20257cb, 32'hb160f01c, 32'hb2cf7b2f, 32'h476b03e4, 32'h3c655a79, 32'hfbd25111, 32'h635e6090, 32'h93262b89, 32'h84182f13, 32'hccf1775a, 32'h90e1b79f, 32'ha1089ccc, 32'h6e470ab0, 32'hcdc0bca5, 32'h6e883bc3, 32'h70f5dbdf, 32'h7c2785be, 32'h445002d6, 32'hb58371d7, 32'hc332a296, 32'hb820c082, 32'hdf072b73, 32'h4f2742fb, 32'hfae1a83b, 32'hae8b29ba, 32'h4295c446, 32'h29305a78, 32'h911df72d, 32'h956a824c, 32'h6dbf1beb, 32'hb2d5f644, 32'h96c205e0, 32'ha3259f34, 32'h9f40d4bb, 32'h79d7725f, 32'h190661df, 32'h8c633866, 32'h52872ca8, 32'hc84fa3a6, 32'h93c5d7f6, 32'habe66206, 32'h21ef7fff, 32'hec9df3c8, 32'h9ff00bf9, 32'he70ce981, 32'hffa51997, 32'h20ee1a6e, 32'h1389dbc8, 32'h26be7ab7, 32'hb4710768, 32'h6334eefb, 32'h4cebdc67, 32'hbe277a5e, 32'h7ec3dda6, 32'h16f3aeb7, 32'hc90a91b7, 32'hcf2c8f44, 32'h59e44c20, 32'hfa75baa0, 32'hf476e58e, 32'h8c53ebac, 32'hba7c2f70, 32'ha14047c1, 32'hc9bd6a16, 32'h255c0cfa, 32'h8e71c77e, 32'hd0288787, 32'h3ab00297, 32'hf5c65823, 32'h19164704, 32'h1164311c, 32'h1d5e1c49, 32'h6571a725, 32'h8277dd5c, 32'h88b8a3a2, 32'h2ab2ef23, 32'hdc778c57, 32'he5b8bd63, 32'h7a836432, 32'h463193cb, 32'h544f4bf2, 32'he5bb8851, 32'h3579d44a, 32'ha7adc50f, 32'h62d3ebfc, 32'h7aa4c035, 32'h37ad2b06, 32'hb5d8b84a, 32'he198f92e, 32'ha71b1ce5, 32'h8be33bc4, 32'hfc30bc20, 32'h4cae94a7, 32'h1b68b5b5, 32'h85a59999, 32'h52cc7af9, 32'h56b9e109, 32'h9dbb2da7, 32'hb89b03e5, 32'ha7f86097, 32'h54e3fae5, 32'hf0e63807, 32'hf1207944, 32'heff5170f, 32'h540cf995, 32'h9457f4b5, 32'h7a1ab137, 32'hf35ec6c3, 32'hf7571b8e, 32'h843c5c71, 32'h325d9488, 32'haeda6bdc, 32'h1e3ee86e, 32'h7fa1d45a, 32'h4d994051, 32'h49a42e30, 32'hfd92707b, 32'hd525b00f, 32'h1dea08b3, 32'hf06fceb4, 32'h556c2a34, 32'hdbfbbb6a, 32'h8054f6f4, 32'h35ed79d8, 32'h4fb90ef1, 32'hb1e13581, 32'h5d320fe4, 32'h32fd0e91, 32'h5627c1ef, 32'h251af3e7, 32'h252a4f76, 32'h2ce56e0d, 32'h95be8f60, 32'hde827528, 32'h1684a374, 32'hd16fb6d9, 32'hb0b7164c, 32'he7664b63, 32'h95e0c963, 32'hb6137db9, 32'h8ce011de, 32'h896315e5, 32'h53a48fee, 32'hf8c4d90d, 32'h4e599a05, 32'hf5435018, 32'h240c5779, 32'h45e0e11d, 32'h985b4ad1, 32'h29e01609, 32'ha607703e, 32'h24f0cb8a, 32'hb1508d73, 32'he6f998b0, 32'hf6c7045b, 32'h71825c6b, 32'h551de9f3, 32'ha16a45bf, 32'he2e0ee2e, 32'hc7e29cf8, 32'h103f76a1, 32'hadb08ecd, 32'h3c18f311, 32'h67729d77, 32'h16a69bfc, 32'hfb89dbe9, 32'h743b54d6, 32'habf9ed46, 32'h5ac98f11, 32'ha1c93ade, 32'hdb0d9837, 32'hae8285d6, 32'h6fb11540, 32'h34fa9fd4, 32'h5aa4a495, 32'hb3b226a3, 32'h3841bdf0, 32'hce0c1dd4, 32'h2c8db8cb, 32'h8323137d, 32'h94d2f788, 32'h40975434, 32'hb96c2d6c, 32'h5efebaf9, 32'hac187616, 32'h478d1530, 32'h4b8bf7e6, 32'hfccd7654, 32'hbb57bd02, 32'ha61abfe9, 32'hac3de853, 32'h56c1cb7b, 32'hf233217f, 32'h4378e685, 32'hc41bddad, 32'h42d028a8, 32'h499f723f, 32'hba93d6d5, 32'h6da9dd0c, 32'he8b461c0, 32'h25b2c5df, 32'h29435464, 32'h2e57e9f6, 32'h1975717d, 32'he2f9d6f7, 32'ha14d20cf, 32'h1a6da9a9, 32'h5ab60804, 32'hd28d0d58, 32'h7e0d5ca1, 32'h4de4f1ea, 32'ha496b5d5, 32'h17d5a39e, 32'h97bba6f9, 32'h4e365c95, 32'h4bdef53f, 32'hcfeb2970, 32'h23f72fd0, 32'h90136635, 32'h8bb1c9dc, 32'hfcb30098, 32'hefdd03b7, 32'h6dd20baf, 32'ha49c770c, 32'hd0c51c89, 32'h55cb2153, 32'he8b335d3, 32'hdf14d3b5, 32'hff7e0293, 32'h56c14001, 32'hfd879862, 32'hc04ce73d, 32'hbd8adbc6, 32'heccf96f8, 32'h947a9311, 32'h536de880, 32'h6f26aaed, 32'h5826d90a, 32'h20bfa689, 32'h1bdae9f4, 32'h6ee25547, 32'h2a974596, 32'h8ea110c4, 32'h3f915c54, 32'h1a8464c1, 32'hacebf11d, 32'hbc8ba464, 32'hf14ae7f1, 32'hae2b26a4, 32'h73f9dc1e, 32'hf077d5b8, 32'h82b3a42c, 32'he218d035, 32'ha96782ec, 32'h6463d592, 32'hd8d20bc3, 32'he03b0409, 32'hd204cb34, 32'h90a3ff8a, 32'hc8ffe85e, 32'hfab0f8ac, 32'h60110331, 32'hd2177893, 32'h12c8107b, 32'h48867812, 32'hc11e717d, 32'h7ed4f4ad, 32'h9c5373e5, 32'h94239bad, 32'h6ef4a13e, 32'h4c49ec71, 32'hf67ecd01, 32'hbd9b4d76, 32'h92824db2, 32'h4a4eabe2, 32'ha55ae1bc, 32'hc8d4ebef, 32'h95410b28, 32'h9b6fa954, 32'habdf3d9e, 32'h8dcdf6d4, 32'hd330c61c, 32'ha4b942f8, 32'h71e87285, 32'hb8b42029, 32'h97c69546, 32'h342a64a4, 32'hd4d93d52, 32'h190526df, 32'hed6eebe1, 32'h69665300, 32'h3f447cce, 32'h356f1e4b, 32'ha4529da3, 32'h7fea0639, 32'hc80c0640, 32'h80364678, 32'h7ccf8254, 32'hae0e6ba5, 32'hcd21c3b2, 32'hfb47a708, 32'h7fe76985, 32'ha0581196, 32'h7347e518, 32'hf30d9efd, 32'hd1c48596, 32'h137f1a57, 32'h2c2ba353, 32'h237df272, 32'h6d81c324, 32'h3d42353d, 32'hdac13cf9, 32'h7eeafe54, 32'h99bb86db, 32'h3e74432b, 32'h344b71a1, 32'h96151426, 32'h66304acd, 32'h762c8204, 32'h7618c9f7, 32'hf20d7db0, 32'hb8f5baac, 32'hb3d8f7bf, 32'hfbcb74a3, 32'he980a384, 32'hd008950c, 32'h4498cf51, 32'hdbd95c46, 32'hf0803639, 32'ha4a77465, 32'haa6e565e, 32'h7f40f29b, 32'h8fb93bfe, 32'h2d57bae1, 32'hb386be4c, 32'h2fc584db, 32'hd66cabda, 32'h412e6aa9, 32'h747071c9, 32'h8295c9ba, 32'hd98fd031, 32'hd4055d14, 32'h990ac741, 32'ha19215b3, 32'h5ca1a729, 32'h1c78c59c, 32'h2f42142b, 32'h3a146f38, 32'h1aa28216, 32'hf769f149, 32'h344204b7, 32'hf2713770, 32'h6e1886e9, 32'hc6d0aeca, 32'h4d04092f, 32'hdf650360, 32'h96d425da, 32'hcf2846a8, 32'h3c30cc0c, 32'h177083c1, 32'h9a7984d6, 32'ha20e42ad, 32'h571238f6, 32'hf6e615dd, 32'h8a602807, 32'hc8bbecda, 32'h75e4f5fd, 32'h2019f9f9, 32'h51604ee9, 32'he18a4005, 32'hf5f71dc6, 32'hc212485c, 32'h73dd3b42, 32'hb302d7fb, 32'h57c97664, 32'h54623b25, 32'ha9c9b07a, 32'h8c1be2b0, 32'ha6b5fb16, 32'h17163f00, 32'h74e3819e, 32'hc1e681b2, 32'h21675aa3, 32'h5d5da4e6, 32'h86eb3630, 32'hdcf410b0, 32'h49a44633, 32'hc269e9c0, 32'h917a5202, 32'h46c7a000, 32'h19895c50, 32'hdc58680d, 32'h45acc069, 32'hb2535a08, 32'h7343133d, 32'h6a883aec, 32'h8182f776, 32'h28a95d01, 32'h30edefd6, 32'h5144fbca, 32'hb1618843, 32'h3d9ef2ca, 32'h617d6418, 32'h46434a0c, 32'h8e4b8cf5, 32'h4ce274bb, 32'h813c902f, 32'h2fe5c25e, 32'hd02764cd, 32'h52e6eaa9, 32'h74c99eea, 32'hbca42c82, 32'hb3777d1f, 32'hee2c450b, 32'h59c584a6, 32'he37afb43, 32'ha807d56b, 32'hd6873020, 32'hc002034a, 32'h838c0934, 32'h6f46f4ab, 32'habc177c0, 32'h533f0918, 32'he81b94c9, 32'hb9b99b54, 32'hd42bf77a, 32'h109a1081, 32'h96bd02cf, 32'h24fe5397, 32'h531becdf, 32'h8783cea5, 32'h8718bf96, 32'h9bc91ae9, 32'h1131bf73, 32'h5cd97f31, 32'h9fade8ad, 32'h8805bad9, 32'hacc82cbb, 32'h116953d8, 32'h7a70e045, 32'h3c69103c, 32'h6abefdd8, 32'h28ad2917, 32'h7cf2d9d1, 32'hc407a241, 32'ha5e8dfdb, 32'hb0d25a2e, 32'h8eb354b8, 32'h147bc2d2, 32'h3c33e1f2, 32'h90c7282b, 32'h6e4f74d8, 32'h8ba6ca7b, 32'hc3ddbed3, 32'h66fdde7e, 32'h3d64a969, 32'h1730d99f, 32'h51dfb083, 32'h17067aa9, 32'h5651ca3c, 32'hbfdd613a, 32'haf285aef, 32'hffa9ed92, 32'hf1cc7f6f, 32'h876a5b16, 32'hbbfb2b6b, 32'h79b4ab03, 32'hecc9f2a2, 32'h8eb63309, 32'h6dc91900, 32'he6d542ce, 32'hbf791827, 32'ha1918970, 32'h333828b6, 32'h112b56b1, 32'he0dca5fd, 32'h925bffc4, 32'h58860809, 32'h99fc4bfe, 32'h406218e4, 32'hc24d14e6, 32'h1b6d3729, 32'h3e870e97, 32'ha86e13df, 32'he89bd896, 32'hc4cfabf5, 32'h68755ce6, 32'h734928aa, 32'h5c8e8010, 32'hf71fd735, 32'hed8b4e52, 32'h7dd969b3, 32'ha6b9bceb, 32'h8d32bf8c, 32'h594676a0, 32'h50621178, 32'hef32c680, 32'h2fdfb11e, 32'h8e751081, 32'hde111a61, 32'had16c940, 32'hc2389c3b, 32'hde1c1aa5, 32'he87f8caf, 32'h242a4477, 32'h9157f463, 32'hd60ac5b7, 32'he2b5e35d, 32'hb65ddfa9, 32'haa0511d6, 32'h521c630e, 32'he498f8ea, 32'haf27de2f, 32'hf95039bc, 32'h652d35d5, 32'h923a5a34, 32'h52035227, 32'h3de7c13f, 32'hdcf96f0e, 32'ha6537c21, 32'h71ee6a7f, 32'hc2c297da, 32'h6fa14588, 32'haf43bee6, 32'h93f93c9a, 32'hfbedea48, 32'h6c2ffa6a, 32'hb7403453, 32'h5c589a0c, 32'h54ffe226, 32'hb88e47ad, 32'hef60578e, 32'hedaaf393, 32'hc9208330, 32'hd8231a78, 32'h332fa37e, 32'h53097101, 32'h3f936455, 32'h1b6fe7b3, 32'h95d23204, 32'he94a62e0, 32'h7b6824c6, 32'h9a706474, 32'h52ce65b3, 32'ha5075090, 32'h17e5e95c, 32'h82973563, 32'ha64a46d0, 32'h4c3b13af, 32'h2bcc6534, 32'h150f2296, 32'ha2c7151e, 32'h165de6e3, 32'h7c9d33b7, 32'h52d74bdc, 32'hafa3f197, 32'h896219a5, 32'h272dd0de, 32'h16411f4d, 32'h1e497009, 32'hee2b42ad, 32'h22020160, 32'h8ca1a4c7, 32'hf720b4f8, 32'h4e6790ce, 32'h9d568cfd, 32'h60d024ce, 32'h36f05531, 32'hc6b86f89, 32'h4fd15420, 32'h139f164a, 32'h55019801, 32'h66ee8eba, 32'h18a2abb0, 32'ha92fcefb, 32'hdddb75e2, 32'h2baba0c9, 32'hc2eb6ade, 32'h8445d72e, 32'h30fc881d, 32'h1a3b2aec, 32'h4593c4eb, 32'h7d68d346, 32'h39d64a6b, 32'h8d00ec0c, 32'h7efe6e60, 32'hae7fb593, 32'h48606478, 32'hc5967d92, 32'hdedb812e, 32'h72f26ad7, 32'h933d824c, 32'h28574ae4, 32'h25270644, 32'hdf3a45ae, 32'h84bded03, 32'h6ecc0146, 32'hccbd772e, 32'h5c46b5d6, 32'h67669f87, 32'h1a0146c7, 32'h4064415a, 32'h7c36d846, 32'h6bfcbe05, 32'h2059e926, 32'h9f0210ad, 32'h476d0efe, 32'hd7615d2e, 32'h94836889, 32'h626bbb04, 32'hf62fd7a5, 32'haca7ce14, 32'hab322cc5, 32'h32d77277, 32'h7e811087, 32'h6723399a, 32'hdb668f55, 32'h466def95, 32'hb3ef7481, 32'h3b6000bd, 32'hc48aa554, 32'he301f5a6, 32'hb8d9f901, 32'h342d71d5, 32'h93344cd4, 32'hb5c0dd79, 32'h36955952, 32'hf8f2d016, 32'he8418e5b, 32'h3305df6b, 32'h9235ac04, 32'h8fa14b5a, 32'h3d3a99c6, 32'h3cfb60bf, 32'h7528685e, 32'hf8fa639a, 32'h51bd8714, 32'h6db49c7d, 32'h8b312c69, 32'heec65457, 32'hdea489db, 32'h9a044fa2, 32'he06093ed, 32'h2960ecb2, 32'h7080a64c, 32'h270e1c54, 32'h5c4e8693, 32'h41c70f32, 32'h4df71c8d, 32'h13da3f6c, 32'h7ee673ec, 32'hbeea63b1, 32'h82fe513a, 32'hd937797e, 32'h11060af1, 32'hc112e2a2, 32'h838e7d02, 32'hdb4e9e19, 32'h8e84b8a1, 32'h8ae13b95, 32'h528d01de, 32'h5425f145, 32'h8d3a3ccd, 32'hf2393f76, 32'h9e803cb0, 32'h33cc5c38, 32'hbfc43eff, 32'h3b0b43d9, 32'h9e983a3e, 32'hcc7d117b, 32'ha3a73882, 32'hfcec8750, 32'hdf75bc31, 32'had1298d2, 32'haf656d16, 32'ha4c976a4, 32'h5d5e3562, 32'h367a4267, 32'hf2f3c53e, 32'h3d59dc9b, 32'hd9d1608e, 32'hd6ac3b25, 32'h5016f4e7, 32'h2cb9572f, 32'hcd9b34ea, 32'haefa6b8a, 32'h3ea12d30, 32'h3b8e95f1, 32'hc1cc6745, 32'ha6ec06a7, 32'h59edcae1, 32'h6ee94a6e, 32'hdc7817e8, 32'he8c91323, 32'hf2598f13, 32'hcd9f7805, 32'h8f7987b0, 32'h2f0c2ae9, 32'h439827ad, 32'h51f90bfd, 32'he2209523, 32'h3c228bad, 32'hec9d3d1f, 32'h151cbdd5, 32'hb3bba2db, 32'h815e9fd2, 32'h69ba7c2e, 32'hbe480b39, 32'h6441773a, 32'h82fbf075, 32'hc0cb9ab1, 32'h6f1a2cf0, 32'hd4258020, 32'hf1cdc683, 32'h3af06f76, 32'hbbd63513, 32'ha0c35a11, 32'h4c7a4b44, 32'h86b71a34, 32'h92e7c715, 32'h44e357a8, 32'hfe50c64e, 32'h187ca2e7, 32'h88cb2b36, 32'he5ac5744, 32'hef068b58, 32'h22709359, 32'h64100167, 32'h3c56ed2e, 32'he19432d8, 32'h28c1d374, 32'hb964f446, 32'hcc708dc3, 32'hb21b7ed1, 32'h199ab159, 32'hb6e53981, 32'hb1e7d8a1, 32'hf0b6cab3, 32'h24cd8b1c, 32'h520bdc1c, 32'hde3fe5b5, 32'h3fea394f, 32'h311611bc, 32'hc77cc7ef, 32'h7cdba692, 32'h5c7b69f5, 32'hcbc2d9c2, 32'h468bec1d, 32'h4e7edd82, 32'h6d0c9a72, 32'hb317ea07, 32'h5ebf1907, 32'hf2461f63, 32'h49cc5cc1, 32'h3dae4aed, 32'h4915da7b, 32'h4ea6e540, 32'hc00706d6, 32'h2559a5d5, 32'hf39b903d, 32'h24cd281f, 32'hef700470, 32'h8b1f79af, 32'h393d386f, 32'he50b4065, 32'h4dca3caa, 32'h549680e1, 32'h9a1bc2be, 32'h345d0623, 32'h3797e56a, 32'he5c61826, 32'h3c38c114, 32'h1468334d, 32'he4e8b9a0, 32'h2a3f8c7c, 32'h9a7871f8, 32'h580a8eb4, 32'h3d8083e6, 32'h8a5ea82a, 32'hff503535, 32'hc57b13f5, 32'h9c5f2fd7, 32'he66c21f2, 32'h1c11e008, 32'h11c2f684, 32'h9962263f, 32'h6c54f489, 32'h9b9adda8, 32'h66d4bb47, 32'he081c615, 32'hcfb7dffb, 32'heec50d32, 32'h87c08fc8, 32'hb028fcde, 32'hac7964fa, 32'h16212ecd, 32'h5e6e16fa, 32'ha3072160, 32'h40b21bc4, 32'h6b3fe4d2, 32'hf7f05140, 32'h66238025, 32'h886e2b4f, 32'hbfbeb6c5, 32'h83066f8e, 32'h98b783b8, 32'h197faab9, 32'h5176e166, 32'h852b8eb6, 32'h5b5db942, 32'h904186a7, 32'h242287cd, 32'h8f057bf2, 32'hb6bd319b, 32'h1911110a, 32'h46402764, 32'hb4926d1c, 32'h6de05d3b, 32'h94e682e9, 32'hcecacc70, 32'h77b4a8e2, 32'h43d898fc, 32'hcaad4c60, 32'h3d9ca43a, 32'h117d8f0f, 32'h4278877b, 32'hba4d2953, 32'h23b6ed70, 32'h6d6ad440, 32'hf72d8fcf, 32'h5e213226, 32'h90a550cb, 32'h153459ec, 32'h6c60d123, 32'hc560d750, 32'ha2f515a2, 32'h2a6b19c4, 32'h5cb9cd18, 32'hb6d62493, 32'h23defb83, 32'h936afb21, 32'h8f1e2552, 32'ha5cd9a2a, 32'haca573e2, 32'ha958f43f, 32'h59b6cfab, 32'hfd513773, 32'h99acadba, 32'h5b953d39, 32'h560e0ada, 32'ha28d4308, 32'h4bf13d43, 32'h59d23e30, 32'h858dca51, 32'hfb774f64, 32'hf948f26f, 32'h91de779e, 32'hf839e403, 32'h43652fe4, 32'h386f39a3, 32'hce6fb2ca, 32'h3ded16e6, 32'hf69762f1, 32'hab0fd05e, 32'hf48079f0, 32'hb008aee8, 32'hdcb677b3, 32'hb461bafa, 32'h3593cf4d, 32'h273c85ee, 32'h10a1b293, 32'h85f94600, 32'hbf04e979, 32'he41dc0b3, 32'hf1408d5d, 32'h591392ca, 32'hda1f7c2e, 32'h6748c520, 32'hfe6077d2, 32'hecf64f09, 32'hf080a2ba, 32'h3562f57a, 32'hb1a40675, 32'h112ba547, 32'hd958c712, 32'h294cfd3e, 32'h8b65e24c, 32'h69aa94c5, 32'hdc5a3db5, 32'hdabe235d, 32'h883c752e, 32'h4e17dc99, 32'hb87f25dc, 32'h5185a9b9, 32'h4dbb462f, 32'h12c0de1e, 32'h95e10359, 32'h863202ea, 32'hfa3572f0, 32'hc8511eba, 32'haf9fab40, 32'h2a4a3e3d, 32'hd399459b, 32'h9c994bc3, 32'h3a523590, 32'h575337d4, 32'h6cf7e8a6, 32'hd6c49fb8, 32'h5c79a9d3, 32'hf571d7de, 32'h4439ab7c, 32'hf64d9738, 32'h299c837b, 32'hc7e4da26, 32'h791b26e1, 32'h8c33fad5, 32'h2c2fa1f0, 32'h52247275, 32'hfc4c94e6, 32'hf7a52675, 32'h2ee54511, 32'hf46d1a94, 32'hb540d4dc, 32'hfd60cf64, 32'h15bca5f1, 32'hf994a305, 32'h10a81683, 32'h9c398324, 32'he3a3d95c, 32'hfd012969, 32'he273bc0a, 32'h2aaeb641, 32'h58d55b3f, 32'hab0c1958, 32'h750583aa, 32'h2d7185f2, 32'h47e28e45, 32'hb1f80c78, 32'hfd6c6c18, 32'h46ad9f5c, 32'h82cf2a52, 32'h9329aaa2, 32'hcf552f5a, 32'hbb6e50fe, 32'hfcbc9302, 32'h967f0c6f, 32'h3e19211e, 32'h34f691d7, 32'h2ade8ae2, 32'ha93c15e9, 32'h629b6c9f, 32'h8e2ec471, 32'ha3b69bbe, 32'h48893088, 32'h58adc8c3, 32'h594343cb, 32'hf60eccae, 32'h2859c14f, 32'h64846ce3, 32'h86eb5cc6, 32'h44ed59c1, 32'h680a7634, 32'h5f7186df, 32'h7ff86e9f, 32'h50b88a8a, 32'h5ce2914e, 32'h3d2c336e, 32'hf179c4f9, 32'h9ce74f36, 32'h31ce50ba, 32'hd2e86169, 32'h8bea7536, 32'h52ea8060, 32'ha7951ef6, 32'h9fee735d, 32'h73c0fbbf, 32'h5b5b3277, 32'h9a1c38d0, 32'h95fd209c, 32'h899468dc, 32'h359ed1a5, 32'h5f318e21, 32'h97b59784, 32'he35d3395, 32'h4122ec79, 32'ha8d733cc, 32'he9cb2751, 32'ha611e007, 32'h430fea49, 32'hd37ae3f8, 32'hebfefb9f, 32'h4e5c3311, 32'hff76850e, 32'hd3d14e55, 32'h89a9cd92, 32'h91109f0b, 32'he2679372, 32'h15d3d9cd, 32'h307c2c7d, 32'h7ef5e322, 32'h2677a8d1, 32'he32f3de7, 32'hd4caebdb, 32'h76991d43, 32'h9bbb4acd, 32'hcc3ae690, 32'h96fdebd1, 32'h5cc794d8, 32'h571518fb, 32'hc6fc62e1, 32'h457cc1ef, 32'hc7c3c151, 32'h13d1820f, 32'hce27b3ee, 32'h4b090234, 32'h9c8a6425, 32'h7f481ce2, 32'h59ec1a16, 32'h26336805, 32'hb0b2688b, 32'h10c145e8, 32'h2d69adc2, 32'hfb2333cb, 32'h69ea7ea7, 32'hf85e4bdf, 32'hd0b8528c, 32'h2ad67b36, 32'hd33f12b3, 32'h7afc630c, 32'h279a66cb, 32'h974a1cc2, 32'hd996c27e, 32'hf7baefa4, 32'h2990e000, 32'hd837758e, 32'hd8b66974, 32'hca426cd3, 32'ha3abf416, 32'ha554fd7a, 32'hb5f50c7b, 32'h4f2de639, 32'h4884fb83, 32'he2cbfe3a, 32'h29f21e27, 32'hc6c83b4d, 32'h513b945e, 32'h27a63ca0, 32'h363f1751, 32'hd3648125, 32'hea65c32a, 32'hba172c72, 32'h1bf653a8, 32'h4b06b274, 32'hb60f6503, 32'hb980d052, 32'h1a63bf5c, 32'hc9b1d8e9, 32'he4408f65, 32'hdcbd92ea, 32'h97a4423c, 32'he51d7f2a, 32'hd3c8f1d9, 32'h9e262312, 32'hca7c0e7a, 32'ha1c536ed, 32'hff9894c6, 32'h735acd9d, 32'hbfccde57, 32'h392fc2d5, 32'h267f2e6f, 32'h6b7c3a7b, 32'h812a2f5d, 32'h509d180a, 32'h6afd4af0, 32'h754f74d2, 32'h50b23297, 32'h43a67b45, 32'h6d90b719, 32'h52cebe8a, 32'hbc9321d3, 32'h2d4da0ec, 32'h2ff241b0, 32'h435cc2ac, 32'h40672438, 32'h5bdd9f49, 32'h33b230ab, 32'h575683b0, 32'hb3694cb2, 32'h3c00d57e, 32'hbadd8e90, 32'hac0a038e, 32'h33400cd5, 32'hbaba9d77, 32'h6d5ae0da, 32'hf06935a0, 32'hd6f63862, 32'h50253ab9, 32'h55ac0a60, 32'h7e5da2ff, 32'h48ccd7f9, 32'h33af32bc, 32'h86a391cb, 32'h838d6cf4, 32'h7012150c, 32'hccef3c3a, 32'h87394e8b, 32'hd4b84350, 32'h71796b82, 32'hb881b7f5, 32'h2a02cc83, 32'hf049dc88, 32'h92dc603c, 32'h9078d7d2, 32'h332e9a5e, 32'h3f138132, 32'h51d7853e, 32'h4e9dbed2, 32'h7f892065, 32'hbe99d6bc, 32'hcdd58a67, 32'h50b6e18d, 32'h2a30d831, 32'h24f1a992, 32'hf3f57d0f, 32'h2c0dd3e5, 32'h605f91d8, 32'h5b1461f2, 32'hbbf7909e, 32'h683c2c7e, 32'hfb3326e1, 32'h48b1d545, 32'hea47e2d4, 32'h4fb0724d, 32'he351c2d7, 32'h1936861a, 32'h9d1b0499, 32'hb1b97596, 32'h5f46ef4c, 32'hb412af93, 32'h82f2f07d, 32'hcd30d0b9, 32'h53785c17, 32'hcda1cd6a, 32'hbf51394c, 32'h4d2e815e, 32'h8800c303, 32'h133f507e, 32'h112613d9, 32'h3c018f65, 32'h3650cdf9, 32'h417b961d, 32'h4756bdc7, 32'h85aa2fa3, 32'h2f387b70, 32'hca632445, 32'hb19c53e7, 32'hc658734d, 32'hc710bd7c, 32'h9635d850, 32'hf0c43eaf, 32'h124bca3d, 32'h895cc30d, 32'h691c34e0, 32'h40917324, 32'h5bd24da3, 32'hd2b5b65f, 32'h7210e7f0, 32'h6f6fbe92, 32'hfdbd8473, 32'h37c0e6d8, 32'h42c08dbc, 32'h6793edd3, 32'he5057495, 32'h2a2cf372, 32'h2a4dbd09, 32'h997a532b, 32'he9475ac3, 32'hda864019, 32'h45822281, 32'hd42944e9, 32'h6996315d, 32'h8ecff4ae, 32'hce4b08d2, 32'h101879fa, 32'hfe68abaa, 32'h44f5d974, 32'hb4dd672d, 32'h20ee8039, 32'he1003cb5, 32'h38469d8c, 32'h970da436, 32'h401fb8cd, 32'h6ba6064b, 32'h4e85f35d, 32'h1d6d22c3, 32'h1907ccae, 32'hb169e3f3, 32'hc1de3831, 32'hb8908b87, 32'hc2b4fc88, 32'hb949dc65, 32'h896cfdb6, 32'h856f29af, 32'h3232f1e1, 32'h9a4aa2fe, 32'h36849a73, 32'hf72458a3, 32'h227ed38e, 32'h20341032, 32'heeed5495, 32'h2eb57161, 32'heeddaed8, 32'h47ca39bd, 32'hf72d30c6, 32'hde6bcaef, 32'h1d8b744c, 32'h41b4d824, 32'h911df5d9, 32'h59c9f76e, 32'h74e57fef, 32'ha4ad792a, 32'h863bd425, 32'hf0090a14, 32'h67b979fc, 32'hf11aab78, 32'ha897b036, 32'h18d14a88, 32'h477f1f6d, 32'h9445d73a, 32'hc54273d4, 32'haeebfa18, 32'he1e785b1, 32'h457098a3, 32'h45036120, 32'h984fbde0, 32'h8e94884f, 32'h6728b5b8, 32'hb6ec3b30, 32'hb130b5e8, 32'h229838b7, 32'h558b6a44, 32'he87a8c43, 32'hbd98ba4b, 32'h831e315b, 32'hab3ee8b4, 32'h6bef7ef5, 32'h2b8df617, 32'h495eff10, 32'hbb48ff10, 32'h6b735dcc, 32'hb75cf8ae, 32'hd546fb79, 32'h7555aa48, 32'h9ee8cbc4, 32'ha031a515, 32'h952bf2dc, 32'habf75cf8, 32'he204bd36, 32'h5685cf78, 32'he40fe5e5, 32'h5e76eca0, 32'hc93b8877, 32'he7f3e69f, 32'h75f09c1f, 32'h6e87df6f, 32'h673931af, 32'hdfbff7f1, 32'hf721eb94, 32'hb6659723, 32'h4a2fbe66, 32'h43626bf5, 32'h32b826f7, 32'hbce098bb, 32'h7a4cbfaa, 32'h6619310d, 32'hf6ebe0d4, 32'h52a176e7, 32'hbe009b78, 32'hbab6f461, 32'he4045205, 32'h9235f613, 32'hab6b7947, 32'ha032d713, 32'hbfb66893, 32'h9b7925a2, 32'ha470a9e1, 32'haeb5c84f, 32'h40cce4bd, 32'h342f4c01, 32'hba82b33a, 32'h3921c0bb, 32'ha960161e, 32'h28437450, 32'h2413c258, 32'h364c4e99, 32'h85f4808b, 32'h1a347251, 32'h46a0a714, 32'he6e05f75, 32'h11437e31, 32'he88d3da1, 32'had7b51c3, 32'hb4816e9b, 32'h99a0e7b7, 32'hda1c7fc9, 32'hc5bbfe7d, 32'hcf49ab14, 32'hd706f6ef, 32'ha44af607, 32'hc8be6587, 32'hfa049ffc, 32'h7fc70226, 32'h44ca6630, 32'h3e153152, 32'ha1a3b986, 32'hdf7dfdfb, 32'h8641503e, 32'h1eef1d83, 32'h2646935c, 32'ha9b86b96, 32'ha7cef756, 32'hc40efd04, 32'h288558cd, 32'h57b2f750, 32'hefde842a, 32'hc77dd5a9, 32'ha54bed54, 32'hc42a6a9c, 32'hc58d8a5e, 32'h8cae786a, 32'h7bbbecff, 32'h3b2400c7, 32'hbfd8b177, 32'h1a183474, 32'h98a3c82a, 32'hcd93dd35, 32'h1e948677, 32'h4005a4e2, 32'h25f3ca55, 32'h5836a593, 32'hfa214c94, 32'h102d858e, 32'h15473846, 32'h1285fb0e, 32'hb50056e8, 32'h690efef1, 32'hdb5a5ed2, 32'h24fa4e36, 32'h70ee9c57, 32'hc50017e6, 32'hd008ddd5, 32'h8b27e002, 32'h25fb95ac, 32'he4cba449, 32'ha515e03d, 32'h26a63fa5, 32'h2043d707, 32'hf94790d4, 32'h5e37d4f0, 32'h9b230b4f, 32'h661f8015, 32'h97fb604a, 32'hecf7779b, 32'h6b0e7498, 32'h843a08c8, 32'ha990cbee, 32'h8ecacb69, 32'h914e70c2, 32'h9fa61503, 32'he300406e, 32'h4e1003d9, 32'h46ef1dca, 32'h22d9d1cc, 32'hc8fc018c, 32'h55a104a4, 32'he4dd7edf, 32'hb657b76f, 32'he052a9d1, 32'hbb11faab, 32'h1d971f95, 32'h156ead46, 32'h18de64cb, 32'hc5e37fa8, 32'h4662c6e2, 32'hcedbe7e9, 32'h5b6be357, 32'hcf355857, 32'h73845657, 32'h1192dabc, 32'h51266d83, 32'hedaab686, 32'h551795c5, 32'h59aafff7, 32'hdf38060f, 32'hc37129f5, 32'ha0b0985d, 32'h8548612f, 32'he878479c, 32'h826a8a4d, 32'h2d53c5ae, 32'hd327cadd, 32'h5d32387a, 32'hf043f80d, 32'hc222e7c8, 32'h6965a055, 32'h6b73a4ec, 32'hce723be8, 32'hf984e8e7, 32'hdf88e157, 32'h77b95e0c, 32'h4cbd9e00, 32'h274032cf, 32'h91611bb0, 32'hd87a1c76, 32'hc3042730, 32'h501fbc8b, 32'hbb8c0f8f, 32'h77f34bed, 32'h2f79de15, 32'h6a18f6e8, 32'h59ad3e7a, 32'h273151cc, 32'h6303b0e7, 32'h9353e463, 32'hc37a18b2, 32'he631d0a1, 32'h99f93772, 32'h67560986, 32'ha0dc579e, 32'h56a22c44, 32'h11a1831e, 32'h1bbc40d6, 32'hbd3cc851, 32'hc287e289, 32'hb694ec9a, 32'h2dd27ce9, 32'h9af2c3c3, 32'hf69630b7, 32'haf280480, 32'h74434031, 32'h5f7565b8, 32'h797f15e2, 32'h6fa827cc, 32'h9abd3c02, 32'ha9e2808b, 32'ha9c15c81, 32'hff11b217, 32'h746d6071, 32'h9a8834bb, 32'h6481e772, 32'hc44e2128, 32'h7d4c6704, 32'h733a91bc, 32'h8e1ce971, 32'h436268f1, 32'h1353124c, 32'hff354a0d, 32'h2407d0e4, 32'h46182442, 32'h63aebb25, 32'h942ef980, 32'hdd9efb79, 32'hdda054ce, 32'h24189267, 32'h7d17395f, 32'h1971f22d, 32'h19c33971, 32'h9a20f0ee, 32'hfb250d6a, 32'he02e0436, 32'he25aa854, 32'h27cbfe0c, 32'h98e46504, 32'h131f7f92, 32'hdb708179, 32'h77e8be0b, 32'h712516ba, 32'h46437f3f, 32'hb44a1b7e, 32'hc965cbc3, 32'hbee3b84c, 32'h96d5c84a, 32'h35f7ccd6, 32'h7f51d8e0, 32'h4302d880, 32'h876edf23, 32'he2963a8d, 32'hff2f231a, 32'h40bbffb9, 32'h37e64adb, 32'h614257b9, 32'ha17e5754, 32'he9b37f59, 32'hcd9890e7, 32'hb8fedc72, 32'h80008b1a, 32'hb5fa80ed, 32'hc4e9f9f0, 32'hd39f9977, 32'hd535eb8b, 32'h39f5307f, 32'hc00b5aaa, 32'hbfe403d1, 32'hed0d6c60, 32'haa0178f4, 32'h3b0bd9b5, 32'h6ce0a73a, 32'hcf36668b, 32'h23d6ba51, 32'hfb79fa69, 32'h4db9d1f1, 32'ha3bd73d7, 32'hfcb07110, 32'h58f71a90, 32'h5488daba, 32'hac6fe2fa, 32'h8022305b, 32'hf6863a79, 32'hd7cb85d0, 32'hfc98a59b, 32'h2f0534de, 32'h34afd968, 32'h66adca1d, 32'h65272c39, 32'h22d815e4, 32'h9bf8f7d3, 32'h4a512deb, 32'h21e35c1d, 32'h4f372407, 32'h714c9106, 32'h2ea839c2, 32'hb388e643, 32'h262ef4c7, 32'h525840a4, 32'h32d5d2c6, 32'hf0a29312, 32'hba3196ec, 32'hfa4c7159, 32'hc1629dc8, 32'hfde41258, 32'hfae87051, 32'h9f74f0be, 32'h3c8716d1, 32'hce30d9c4, 32'hccc01157, 32'h4d3fdf48, 32'h97816c3b, 32'he4f9ea4f, 32'h36c03a27, 32'hc6e03466, 32'h9adef997, 32'h9d8e3d30, 32'h7af75766, 32'h8629a590, 32'hfa6df5ac, 32'h6afb055f, 32'hefe3cc73, 32'hf2bed5ac, 32'hc2fdec33, 32'h3e853ab5, 32'h9ddbd992, 32'h9cc52d71, 32'h52a82a63, 32'h29eb5193, 32'h165622db, 32'h57addaa6, 32'h92cf304b, 32'h96a880b3, 32'h606cf49e, 32'h769197cf, 32'h21029f36, 32'h298a4426, 32'h579d5442, 32'h3ef0a30a, 32'hd765f55e, 32'h11dfc3bf, 32'ha6a1f973, 32'hd8b08151, 32'h6937bd7d, 32'h13f99abb, 32'h350662a4, 32'h1ccd183c, 32'h356c6398, 32'hfbc8a667, 32'h6ce0ea70, 32'h1b56c074, 32'h7577975e, 32'h381693d4, 32'h76894406, 32'h6e1512d2, 32'h510bd851, 32'h7dcb8701, 32'h36748d35, 32'h31f76bb9, 32'h72602b94, 32'h96f56738, 32'hf21a6b2d, 32'h28c10f1b, 32'h74e10773, 32'had64b146, 32'h6649cca5, 32'ha38c43ee, 32'h88aa66af, 32'h995fa1f5, 32'hd9660c9f, 32'hd3dee4a8, 32'h3c724c47, 32'h1ebc4f1d, 32'h60a3a7e0, 32'h472a2e11, 32'hb4e5c951, 32'h61302212, 32'hcf5f2abb, 32'h1583c765, 32'hf50e04bb, 32'h5e0d6413, 32'h8300845d, 32'h5125da05, 32'h1d568e59, 32'he9199297, 32'h92e8d880, 32'h1b22ddf3, 32'h43a15294, 32'hfd32e8e8, 32'h7a64f6b2, 32'h90c05244, 32'h6f0a39b0, 32'h9c773fea, 32'he68dfcdd, 32'h26b0ccb3, 32'h2ef42eab, 32'h4fbb5314, 32'hb792b1e6, 32'h4d411f9b, 32'hef23e6ac, 32'hc035b3ff, 32'hb0ab63b3, 32'h2efff576, 32'h2f462279, 32'h8dacb848, 32'h9859b4de, 32'h9c45d971, 32'h44928edf, 32'hd87ff21b, 32'h269b1443, 32'h6dac1191, 32'he5e49802, 32'h1728648d, 32'h6d346403, 32'hec7c16b7, 32'hc02818f5, 32'h82a6ff28, 32'h76c5cc80, 32'hc6cec170, 32'h60c8b455, 32'hed3032a8, 32'hd370e540, 32'h55c38ebc, 32'h29742c41, 32'h627ce300, 32'h40ed025b, 32'hb5b70d8f, 32'hb51b672e, 32'h199c452b};
    
    wire [63:0] bits [N_CORES-1:0];
	wire [63:0] bit_errors_pre[N_CORES-1:0];
	wire [63:0] bit_errors_post[N_CORES-1:0];
	wire [63:0] frames[N_CORES-1:0];
	wire [63:0] frame_errors[N_CORES-1:0];
    
    genvar i;
    
    generate
        for (i=0; i < N_CORES; i=i+1) begin
            sys3 #(
                .RANDOM_64(RANDOM_64[(i+1)*4-1:i*4])
                ) core (
                .clk(clk),
                .rstn(rstn),
                .en(en),
                .probability_in(probability_in),
                .probability_idx(probability_idx),
                //.precode_en(precode_en),
                .n_interleave(n_interleave),
                //.ifec_en(ifec_en),
               .total_bits(bits[i]),
               .total_bit_errors_pre(bit_errors_pre[i]),
               .total_bit_errors_post(bit_errors_post[i]),
               .total_frames(frames[i]),
               .total_frame_errors(frame_errors[i]));
        end
    endgenerate 
    
    
    // below is to sum all bits and bit errors across cores
    wire [63:0] bits_summation [N_CORES-1 : 0];
    wire [63:0] bit_errors_pre_summation [N_CORES-1 : 0];
    wire [63:0] bit_errors_post_summation [N_CORES-1 : 0];
    wire [63:0] frames_summation [N_CORES-1 : 0];
    wire [63:0] frame_errors_summation [N_CORES-1 : 0];
    
    generate
        
        for(i=0; i<N_CORES; i=i+1) begin
        
            if (i == 0) begin
                assign bits_summation[0] = bits[0];
                assign bit_errors_pre_summation[0] = bit_errors_pre[0];
                assign bit_errors_post_summation[0] = bit_errors_post[0];
                assign frames_summation[0] = frames[0];
                assign frame_errors_summation[0] = frame_errors[0];

                
            end else begin
                assign bits_summation[i] = bits_summation[i-1] + bits[i];
                assign bit_errors_pre_summation[i] = bit_errors_pre_summation[i-1] + bit_errors_pre[i];
                assign bit_errors_post_summation[i] = bit_errors_post_summation[i-1] + bit_errors_post[i];
                assign frames_summation[i] = frames_summation[i-1] + frames[i];
                assign frame_errors_summation[i] = frame_errors_summation[i-1] + frame_errors[i];

            end
        end
    endgenerate
    
    assign total_bits = bits_summation[N_CORES-1];
    assign total_bit_errors_pre = bit_errors_pre_summation[N_CORES-1];
    assign total_bit_errors_post = bit_errors_post_summation[N_CORES-1];
    assign total_frames = frames_summation[N_CORES-1];
    assign total_frame_errors = frame_errors_summation[N_CORES-1];
    
endmodule


